// (C) 2001-2012 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// $Id: //acds/rel/12.1/ip/merlin/altera_merlin_router/altera_merlin_router.sv.terp#1 $
// $Revision: #1 $
// $Date: 2012/08/12 $
// $Author: swbranch $

// -------------------------------------------------------
// Merlin Router
//
// Asserts the appropriate one-hot encoded channel based on 
// either (a) the address or (b) the dest id. The DECODER_TYPE
// parameter controls this behaviour. 0 means address decoder,
// 1 means dest id decoder.
//
// In the case of (a), it also sets the destination id.
// -------------------------------------------------------

`timescale 1 ns / 1 ns

module SoC_addr_router_006_default_decode
  #(
     parameter DEFAULT_CHANNEL = 0,
               DEFAULT_DESTID = 1 
   )
  (output [96 - 91 : 0] default_destination_id,
   output [55-1 : 0] default_src_channel
  );

  assign default_destination_id = 
    DEFAULT_DESTID[96 - 91 : 0];
  generate begin : default_decode
    if (DEFAULT_CHANNEL == -1)
      assign default_src_channel = '0;
    else
      assign default_src_channel = 55'b1 << DEFAULT_CHANNEL;
  end
  endgenerate

endmodule


module SoC_addr_router_006
(
    // -------------------
    // Clock & Reset
    // -------------------
    input clk,
    input reset,

    // -------------------
    // Command Sink (Input)
    // -------------------
    input                       sink_valid,
    input  [107-1 : 0]    sink_data,
    input                       sink_startofpacket,
    input                       sink_endofpacket,
    output                      sink_ready,

    // -------------------
    // Command Source (Output)
    // -------------------
    output                          src_valid,
    output reg [107-1    : 0] src_data,
    output reg [55-1 : 0] src_channel,
    output                          src_startofpacket,
    output                          src_endofpacket,
    input                           src_ready
);

    // -------------------------------------------------------
    // Local parameters and variables
    // -------------------------------------------------------
    localparam PKT_ADDR_H = 63;
    localparam PKT_ADDR_L = 36;
    localparam PKT_DEST_ID_H = 96;
    localparam PKT_DEST_ID_L = 91;
    localparam ST_DATA_W = 107;
    localparam ST_CHANNEL_W = 55;
    localparam DECODER_TYPE = 0;

    localparam PKT_TRANS_WRITE = 66;
    localparam PKT_TRANS_READ  = 67;

    localparam PKT_ADDR_W = PKT_ADDR_H-PKT_ADDR_L + 1;
    localparam PKT_DEST_ID_W = PKT_DEST_ID_H-PKT_DEST_ID_L + 1;




    // -------------------------------------------------------
    // Figure out the number of bits to mask off for each slave span
    // during address decoding
    // -------------------------------------------------------
    localparam PAD0 = log2ceil(64'h8000000 - 64'h0);
    localparam PAD1 = log2ceil(64'h8001000 - 64'h8000800);
    localparam PAD2 = log2ceil(64'h8001020 - 64'h8001000);
    localparam PAD3 = log2ceil(64'h8001040 - 64'h8001020);
    localparam PAD4 = log2ceil(64'h8001048 - 64'h8001040);
    localparam PAD5 = log2ceil(64'h800104c - 64'h8001048);
    localparam PAD6 = log2ceil(64'h8001050 - 64'h800104c);
    localparam PAD7 = log2ceil(64'h8001054 - 64'h8001050);
    localparam PAD8 = log2ceil(64'h8001058 - 64'h8001054);
    localparam PAD9 = log2ceil(64'h8001080 - 64'h8001060);
    localparam PAD10 = log2ceil(64'h80010a0 - 64'h8001080);
    localparam PAD11 = log2ceil(64'h80010c0 - 64'h80010a0);
    localparam PAD12 = log2ceil(64'h8001c00 - 64'h8001800);
    // -------------------------------------------------------
    // Work out which address bits are significant based on the
    // address range of the slaves. If the required width is too
    // large or too small, we use the address field width instead.
    // -------------------------------------------------------
    localparam ADDR_RANGE = 64'h8001c00;
    localparam RANGE_ADDR_WIDTH = log2ceil(ADDR_RANGE);
    localparam OPTIMIZED_ADDR_H = (RANGE_ADDR_WIDTH > PKT_ADDR_W) ||
                                  (RANGE_ADDR_WIDTH == 0) ?
                                        PKT_ADDR_H :
                                        PKT_ADDR_L + RANGE_ADDR_WIDTH - 1;
    localparam RG = RANGE_ADDR_WIDTH-1;

      wire [PKT_ADDR_W-1 : 0] address = sink_data[OPTIMIZED_ADDR_H : PKT_ADDR_L];

    // -------------------------------------------------------
    // Pass almost everything through, untouched
    // -------------------------------------------------------
    assign sink_ready        = src_ready;
    assign src_valid         = sink_valid;
    assign src_startofpacket = sink_startofpacket;
    assign src_endofpacket   = sink_endofpacket;

    wire [PKT_DEST_ID_W-1:0] default_destid;
    wire [55-1 : 0] default_src_channel;




    SoC_addr_router_006_default_decode the_default_decode(
      .default_destination_id (default_destid),
      .default_src_channel (default_src_channel)
    );

    always @* begin
        src_data    = sink_data;
        src_channel = default_src_channel;

        src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = default_destid;
        // --------------------------------------------------
        // Address Decoder
        // Sets the channel and destination ID based on the address
        // --------------------------------------------------

        // ( 0x0 .. 0x8000000 )
        if ( {address[RG:PAD0],{PAD0{1'b0}}} == 28'h0 ) begin
            src_channel = 55'b0000000000001;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 1;
        end

        // ( 0x8000800 .. 0x8001000 )
        if ( {address[RG:PAD1],{PAD1{1'b0}}} == 28'h8000800 ) begin
            src_channel = 55'b0000000100000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 33;
        end

        // ( 0x8001000 .. 0x8001020 )
        if ( {address[RG:PAD2],{PAD2{1'b0}}} == 28'h8001000 ) begin
            src_channel = 55'b1000000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 40;
        end

        // ( 0x8001020 .. 0x8001040 )
        if ( {address[RG:PAD3],{PAD3{1'b0}}} == 28'h8001020 ) begin
            src_channel = 55'b0000010000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 35;
        end

        // ( 0x8001040 .. 0x8001048 )
        if ( {address[RG:PAD4],{PAD4{1'b0}}} == 28'h8001040 ) begin
            src_channel = 55'b0000001000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 34;
        end

        // ( 0x8001048 .. 0x800104c )
        if ( {address[RG:PAD5],{PAD5{1'b0}}} == 28'h8001048 ) begin
            src_channel = 55'b0100000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 39;
        end

        // ( 0x800104c .. 0x8001050 )
        if ( {address[RG:PAD6],{PAD6{1'b0}}} == 28'h800104c ) begin
            src_channel = 55'b0010000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 38;
        end

        // ( 0x8001050 .. 0x8001054 )
        if ( {address[RG:PAD7],{PAD7{1'b0}}} == 28'h8001050 ) begin
            src_channel = 55'b0001000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 37;
        end

        // ( 0x8001054 .. 0x8001058 )
        if ( {address[RG:PAD8],{PAD8{1'b0}}} == 28'h8001054 ) begin
            src_channel = 55'b0000100000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 36;
        end

        // ( 0x8001060 .. 0x8001080 )
        if ( {address[RG:PAD9],{PAD9{1'b0}}} == 28'h8001060 ) begin
            src_channel = 55'b0000000001000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 9;
        end

        // ( 0x8001080 .. 0x80010a0 )
        if ( {address[RG:PAD10],{PAD10{1'b0}}} == 28'h8001080 ) begin
            src_channel = 55'b0000000000100;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 8;
        end

        // ( 0x80010a0 .. 0x80010c0 )
        if ( {address[RG:PAD11],{PAD11{1'b0}}} == 28'h80010a0 ) begin
            src_channel = 55'b0000000000010;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 5;
        end

        // ( 0x8001800 .. 0x8001c00 )
        if ( {address[RG:PAD12],{PAD12{1'b0}}} == 28'h8001800 ) begin
            src_channel = 55'b0000000010000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 32;
        end

end


    // --------------------------------------------------
    // Ceil(log2()) function
    // --------------------------------------------------
    function integer log2ceil;
        input reg[65:0] val;
        reg [65:0] i;

        begin
            i = 1;
            log2ceil = 0;

            while (i < val) begin
                log2ceil = log2ceil + 1;
                i = i << 1;
            end
        end
    endfunction

endmodule


