// SoC.v

// Generated using ACDS version 12.1 177 at 2023.01.14.09:41:06

`timescale 1 ps / 1 ps
module SoC (
		output wire [12:0] sdram_controller_wire_addr,  // sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,    //                      .ba
		output wire        sdram_controller_wire_cas_n, //                      .cas_n
		output wire        sdram_controller_wire_cke,   //                      .cke
		output wire        sdram_controller_wire_cs_n,  //                      .cs_n
		inout  wire [31:0] sdram_controller_wire_dq,    //                      .dq
		output wire [3:0]  sdram_controller_wire_dqm,   //                      .dqm
		output wire        sdram_controller_wire_ras_n, //                      .ras_n
		output wire        sdram_controller_wire_we_n,  //                      .we_n
		output wire        c0_clk,                      //                    c0.clk
		input  wire        reset_reset_n,               //                 reset.reset_n
		input  wire        clk_clk                      //                   clk.clk
	);

	wire          cpu_2_jtag_debug_module_reset_reset;                                                                // cpu_2:jtag_debug_module_resetrequest -> [id_router_043:reset, jtag_uart_2:rst_n, jtag_uart_2_avalon_jtag_slave_translator:reset, jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_043:reset, rst_controller_003:reset_in1, rst_controller_011:reset_in2, rst_controller_012:reset_in1, rst_controller_015:reset_in3]
	wire          cpu_0_instruction_master_waitrequest;                                                               // cpu_0_instruction_master_translator:av_waitrequest -> cpu_0:i_waitrequest
	wire   [27:0] cpu_0_instruction_master_address;                                                                   // cpu_0:i_address -> cpu_0_instruction_master_translator:av_address
	wire          cpu_0_instruction_master_read;                                                                      // cpu_0:i_read -> cpu_0_instruction_master_translator:av_read
	wire   [31:0] cpu_0_instruction_master_readdata;                                                                  // cpu_0_instruction_master_translator:av_readdata -> cpu_0:i_readdata
	wire          cpu_0_instruction_master_readdatavalid;                                                             // cpu_0_instruction_master_translator:av_readdatavalid -> cpu_0:i_readdatavalid
	wire          cpu_0_data_master_waitrequest;                                                                      // cpu_0_data_master_translator:av_waitrequest -> cpu_0:d_waitrequest
	wire   [31:0] cpu_0_data_master_writedata;                                                                        // cpu_0:d_writedata -> cpu_0_data_master_translator:av_writedata
	wire   [27:0] cpu_0_data_master_address;                                                                          // cpu_0:d_address -> cpu_0_data_master_translator:av_address
	wire          cpu_0_data_master_write;                                                                            // cpu_0:d_write -> cpu_0_data_master_translator:av_write
	wire          cpu_0_data_master_read;                                                                             // cpu_0:d_read -> cpu_0_data_master_translator:av_read
	wire   [31:0] cpu_0_data_master_readdata;                                                                         // cpu_0_data_master_translator:av_readdata -> cpu_0:d_readdata
	wire          cpu_0_data_master_debugaccess;                                                                      // cpu_0:jtag_debug_module_debugaccess_to_roms -> cpu_0_data_master_translator:av_debugaccess
	wire    [3:0] cpu_0_data_master_byteenable;                                                                       // cpu_0:d_byteenable -> cpu_0_data_master_translator:av_byteenable
	wire          cpu_5_data_master_waitrequest;                                                                      // cpu_5_data_master_translator:av_waitrequest -> cpu_5:d_waitrequest
	wire   [31:0] cpu_5_data_master_writedata;                                                                        // cpu_5:d_writedata -> cpu_5_data_master_translator:av_writedata
	wire   [27:0] cpu_5_data_master_address;                                                                          // cpu_5:d_address -> cpu_5_data_master_translator:av_address
	wire          cpu_5_data_master_write;                                                                            // cpu_5:d_write -> cpu_5_data_master_translator:av_write
	wire          cpu_5_data_master_read;                                                                             // cpu_5:d_read -> cpu_5_data_master_translator:av_read
	wire   [31:0] cpu_5_data_master_readdata;                                                                         // cpu_5_data_master_translator:av_readdata -> cpu_5:d_readdata
	wire          cpu_5_data_master_debugaccess;                                                                      // cpu_5:jtag_debug_module_debugaccess_to_roms -> cpu_5_data_master_translator:av_debugaccess
	wire    [3:0] cpu_5_data_master_byteenable;                                                                       // cpu_5:d_byteenable -> cpu_5_data_master_translator:av_byteenable
	wire          cpu_1_instruction_master_waitrequest;                                                               // cpu_1_instruction_master_translator:av_waitrequest -> cpu_1:i_waitrequest
	wire   [27:0] cpu_1_instruction_master_address;                                                                   // cpu_1:i_address -> cpu_1_instruction_master_translator:av_address
	wire          cpu_1_instruction_master_read;                                                                      // cpu_1:i_read -> cpu_1_instruction_master_translator:av_read
	wire   [31:0] cpu_1_instruction_master_readdata;                                                                  // cpu_1_instruction_master_translator:av_readdata -> cpu_1:i_readdata
	wire          cpu_1_instruction_master_readdatavalid;                                                             // cpu_1_instruction_master_translator:av_readdatavalid -> cpu_1:i_readdatavalid
	wire          cpu_1_data_master_waitrequest;                                                                      // cpu_1_data_master_translator:av_waitrequest -> cpu_1:d_waitrequest
	wire   [31:0] cpu_1_data_master_writedata;                                                                        // cpu_1:d_writedata -> cpu_1_data_master_translator:av_writedata
	wire   [27:0] cpu_1_data_master_address;                                                                          // cpu_1:d_address -> cpu_1_data_master_translator:av_address
	wire          cpu_1_data_master_write;                                                                            // cpu_1:d_write -> cpu_1_data_master_translator:av_write
	wire          cpu_1_data_master_read;                                                                             // cpu_1:d_read -> cpu_1_data_master_translator:av_read
	wire   [31:0] cpu_1_data_master_readdata;                                                                         // cpu_1_data_master_translator:av_readdata -> cpu_1:d_readdata
	wire          cpu_1_data_master_debugaccess;                                                                      // cpu_1:jtag_debug_module_debugaccess_to_roms -> cpu_1_data_master_translator:av_debugaccess
	wire    [3:0] cpu_1_data_master_byteenable;                                                                       // cpu_1:d_byteenable -> cpu_1_data_master_translator:av_byteenable
	wire          cpu_2_data_master_waitrequest;                                                                      // cpu_2_data_master_translator:av_waitrequest -> cpu_2:d_waitrequest
	wire   [31:0] cpu_2_data_master_writedata;                                                                        // cpu_2:d_writedata -> cpu_2_data_master_translator:av_writedata
	wire   [27:0] cpu_2_data_master_address;                                                                          // cpu_2:d_address -> cpu_2_data_master_translator:av_address
	wire          cpu_2_data_master_write;                                                                            // cpu_2:d_write -> cpu_2_data_master_translator:av_write
	wire          cpu_2_data_master_read;                                                                             // cpu_2:d_read -> cpu_2_data_master_translator:av_read
	wire   [31:0] cpu_2_data_master_readdata;                                                                         // cpu_2_data_master_translator:av_readdata -> cpu_2:d_readdata
	wire          cpu_2_data_master_debugaccess;                                                                      // cpu_2:jtag_debug_module_debugaccess_to_roms -> cpu_2_data_master_translator:av_debugaccess
	wire    [3:0] cpu_2_data_master_byteenable;                                                                       // cpu_2:d_byteenable -> cpu_2_data_master_translator:av_byteenable
	wire          cpu_3_data_master_waitrequest;                                                                      // cpu_3_data_master_translator:av_waitrequest -> cpu_3:d_waitrequest
	wire   [31:0] cpu_3_data_master_writedata;                                                                        // cpu_3:d_writedata -> cpu_3_data_master_translator:av_writedata
	wire   [27:0] cpu_3_data_master_address;                                                                          // cpu_3:d_address -> cpu_3_data_master_translator:av_address
	wire          cpu_3_data_master_write;                                                                            // cpu_3:d_write -> cpu_3_data_master_translator:av_write
	wire          cpu_3_data_master_read;                                                                             // cpu_3:d_read -> cpu_3_data_master_translator:av_read
	wire   [31:0] cpu_3_data_master_readdata;                                                                         // cpu_3_data_master_translator:av_readdata -> cpu_3:d_readdata
	wire          cpu_3_data_master_debugaccess;                                                                      // cpu_3:jtag_debug_module_debugaccess_to_roms -> cpu_3_data_master_translator:av_debugaccess
	wire    [3:0] cpu_3_data_master_byteenable;                                                                       // cpu_3:d_byteenable -> cpu_3_data_master_translator:av_byteenable
	wire          cpu_2_instruction_master_waitrequest;                                                               // cpu_2_instruction_master_translator:av_waitrequest -> cpu_2:i_waitrequest
	wire   [27:0] cpu_2_instruction_master_address;                                                                   // cpu_2:i_address -> cpu_2_instruction_master_translator:av_address
	wire          cpu_2_instruction_master_read;                                                                      // cpu_2:i_read -> cpu_2_instruction_master_translator:av_read
	wire   [31:0] cpu_2_instruction_master_readdata;                                                                  // cpu_2_instruction_master_translator:av_readdata -> cpu_2:i_readdata
	wire          cpu_2_instruction_master_readdatavalid;                                                             // cpu_2_instruction_master_translator:av_readdatavalid -> cpu_2:i_readdatavalid
	wire          cpu_3_instruction_master_waitrequest;                                                               // cpu_3_instruction_master_translator:av_waitrequest -> cpu_3:i_waitrequest
	wire   [27:0] cpu_3_instruction_master_address;                                                                   // cpu_3:i_address -> cpu_3_instruction_master_translator:av_address
	wire          cpu_3_instruction_master_read;                                                                      // cpu_3:i_read -> cpu_3_instruction_master_translator:av_read
	wire   [31:0] cpu_3_instruction_master_readdata;                                                                  // cpu_3_instruction_master_translator:av_readdata -> cpu_3:i_readdata
	wire          cpu_3_instruction_master_readdatavalid;                                                             // cpu_3_instruction_master_translator:av_readdatavalid -> cpu_3:i_readdatavalid
	wire          cpu_4_data_master_waitrequest;                                                                      // cpu_4_data_master_translator:av_waitrequest -> cpu_4:d_waitrequest
	wire   [31:0] cpu_4_data_master_writedata;                                                                        // cpu_4:d_writedata -> cpu_4_data_master_translator:av_writedata
	wire   [27:0] cpu_4_data_master_address;                                                                          // cpu_4:d_address -> cpu_4_data_master_translator:av_address
	wire          cpu_4_data_master_write;                                                                            // cpu_4:d_write -> cpu_4_data_master_translator:av_write
	wire          cpu_4_data_master_read;                                                                             // cpu_4:d_read -> cpu_4_data_master_translator:av_read
	wire   [31:0] cpu_4_data_master_readdata;                                                                         // cpu_4_data_master_translator:av_readdata -> cpu_4:d_readdata
	wire          cpu_4_data_master_debugaccess;                                                                      // cpu_4:jtag_debug_module_debugaccess_to_roms -> cpu_4_data_master_translator:av_debugaccess
	wire    [3:0] cpu_4_data_master_byteenable;                                                                       // cpu_4:d_byteenable -> cpu_4_data_master_translator:av_byteenable
	wire          cpu_4_instruction_master_waitrequest;                                                               // cpu_4_instruction_master_translator:av_waitrequest -> cpu_4:i_waitrequest
	wire   [27:0] cpu_4_instruction_master_address;                                                                   // cpu_4:i_address -> cpu_4_instruction_master_translator:av_address
	wire          cpu_4_instruction_master_read;                                                                      // cpu_4:i_read -> cpu_4_instruction_master_translator:av_read
	wire   [31:0] cpu_4_instruction_master_readdata;                                                                  // cpu_4_instruction_master_translator:av_readdata -> cpu_4:i_readdata
	wire          cpu_4_instruction_master_readdatavalid;                                                             // cpu_4_instruction_master_translator:av_readdatavalid -> cpu_4:i_readdatavalid
	wire          cpu_5_instruction_master_waitrequest;                                                               // cpu_5_instruction_master_translator:av_waitrequest -> cpu_5:i_waitrequest
	wire   [27:0] cpu_5_instruction_master_address;                                                                   // cpu_5:i_address -> cpu_5_instruction_master_translator:av_address
	wire          cpu_5_instruction_master_read;                                                                      // cpu_5:i_read -> cpu_5_instruction_master_translator:av_read
	wire   [31:0] cpu_5_instruction_master_readdata;                                                                  // cpu_5_instruction_master_translator:av_readdata -> cpu_5:i_readdata
	wire          cpu_5_instruction_master_readdatavalid;                                                             // cpu_5_instruction_master_translator:av_readdatavalid -> cpu_5:i_readdatavalid
	wire   [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_0_jtag_debug_module_translator:av_writedata -> cpu_0:jtag_debug_module_writedata
	wire    [8:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_0_jtag_debug_module_translator:av_address -> cpu_0:jtag_debug_module_address
	wire          cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_0_jtag_debug_module_translator:av_chipselect -> cpu_0:jtag_debug_module_select
	wire          cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_0_jtag_debug_module_translator:av_write -> cpu_0:jtag_debug_module_write
	wire   [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_0:jtag_debug_module_readdata -> cpu_0_jtag_debug_module_translator:av_readdata
	wire          cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_0_jtag_debug_module_translator:av_begintransfer -> cpu_0:jtag_debug_module_begintransfer
	wire          cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_0_jtag_debug_module_translator:av_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire    [3:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_0_jtag_debug_module_translator:av_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest;                                     // sdram_controller:za_waitrequest -> sdram_controller_s1_translator:av_waitrequest
	wire   [31:0] sdram_controller_s1_translator_avalon_anti_slave_0_writedata;                                       // sdram_controller_s1_translator:av_writedata -> sdram_controller:az_data
	wire   [24:0] sdram_controller_s1_translator_avalon_anti_slave_0_address;                                         // sdram_controller_s1_translator:av_address -> sdram_controller:az_addr
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_chipselect;                                      // sdram_controller_s1_translator:av_chipselect -> sdram_controller:az_cs
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_write;                                           // sdram_controller_s1_translator:av_write -> sdram_controller:az_wr_n
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_read;                                            // sdram_controller_s1_translator:av_read -> sdram_controller:az_rd_n
	wire   [31:0] sdram_controller_s1_translator_avalon_anti_slave_0_readdata;                                        // sdram_controller:za_data -> sdram_controller_s1_translator:av_readdata
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid;                                   // sdram_controller:za_valid -> sdram_controller_s1_translator:av_readdatavalid
	wire    [3:0] sdram_controller_s1_translator_avalon_anti_slave_0_byteenable;                                      // sdram_controller_s1_translator:av_byteenable -> sdram_controller:az_be_n
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire    [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                  // timer_0_s1_translator:av_address -> timer_0:address
	wire          timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire          timer_0_s1_translator_avalon_anti_slave_0_write;                                                    // timer_0_s1_translator:av_write -> timer_0:write_n
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire    [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire          fifo_0_stage1_to_2_in_translator_avalon_anti_slave_0_waitrequest;                                   // fifo_0_stage1_to_2:avalonmm_write_slave_waitrequest -> fifo_0_stage1_to_2_in_translator:av_waitrequest
	wire   [31:0] fifo_0_stage1_to_2_in_translator_avalon_anti_slave_0_writedata;                                     // fifo_0_stage1_to_2_in_translator:av_writedata -> fifo_0_stage1_to_2:avalonmm_write_slave_writedata
	wire          fifo_0_stage1_to_2_in_translator_avalon_anti_slave_0_write;                                         // fifo_0_stage1_to_2_in_translator:av_write -> fifo_0_stage1_to_2:avalonmm_write_slave_write
	wire   [31:0] fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_writedata;                                 // fifo_0_stage1_to_2_in_csr_translator:av_writedata -> fifo_0_stage1_to_2:wrclk_control_slave_writedata
	wire    [2:0] fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_address;                                   // fifo_0_stage1_to_2_in_csr_translator:av_address -> fifo_0_stage1_to_2:wrclk_control_slave_address
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_write;                                     // fifo_0_stage1_to_2_in_csr_translator:av_write -> fifo_0_stage1_to_2:wrclk_control_slave_write
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_read;                                      // fifo_0_stage1_to_2_in_csr_translator:av_read -> fifo_0_stage1_to_2:wrclk_control_slave_read
	wire   [31:0] fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_readdata;                                  // fifo_0_stage1_to_2:wrclk_control_slave_readdata -> fifo_0_stage1_to_2_in_csr_translator:av_readdata
	wire          fifo_1_stage1_to_2_in_translator_avalon_anti_slave_0_waitrequest;                                   // fifo_1_stage1_to_2:avalonmm_write_slave_waitrequest -> fifo_1_stage1_to_2_in_translator:av_waitrequest
	wire   [31:0] fifo_1_stage1_to_2_in_translator_avalon_anti_slave_0_writedata;                                     // fifo_1_stage1_to_2_in_translator:av_writedata -> fifo_1_stage1_to_2:avalonmm_write_slave_writedata
	wire          fifo_1_stage1_to_2_in_translator_avalon_anti_slave_0_write;                                         // fifo_1_stage1_to_2_in_translator:av_write -> fifo_1_stage1_to_2:avalonmm_write_slave_write
	wire          fifo_2_stage1_to_2_in_translator_avalon_anti_slave_0_waitrequest;                                   // fifo_2_stage1_to_2:avalonmm_write_slave_waitrequest -> fifo_2_stage1_to_2_in_translator:av_waitrequest
	wire   [31:0] fifo_2_stage1_to_2_in_translator_avalon_anti_slave_0_writedata;                                     // fifo_2_stage1_to_2_in_translator:av_writedata -> fifo_2_stage1_to_2:avalonmm_write_slave_writedata
	wire          fifo_2_stage1_to_2_in_translator_avalon_anti_slave_0_write;                                         // fifo_2_stage1_to_2_in_translator:av_write -> fifo_2_stage1_to_2:avalonmm_write_slave_write
	wire   [31:0] fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_writedata;                                 // fifo_2_stage1_to_2_in_csr_translator:av_writedata -> fifo_2_stage1_to_2:wrclk_control_slave_writedata
	wire    [2:0] fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_address;                                   // fifo_2_stage1_to_2_in_csr_translator:av_address -> fifo_2_stage1_to_2:wrclk_control_slave_address
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_write;                                     // fifo_2_stage1_to_2_in_csr_translator:av_write -> fifo_2_stage1_to_2:wrclk_control_slave_write
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_read;                                      // fifo_2_stage1_to_2_in_csr_translator:av_read -> fifo_2_stage1_to_2:wrclk_control_slave_read
	wire   [31:0] fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_readdata;                                  // fifo_2_stage1_to_2:wrclk_control_slave_readdata -> fifo_2_stage1_to_2_in_csr_translator:av_readdata
	wire   [31:0] fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_writedata;                                 // fifo_1_stage1_to_2_in_csr_translator:av_writedata -> fifo_1_stage1_to_2:wrclk_control_slave_writedata
	wire    [2:0] fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_address;                                   // fifo_1_stage1_to_2_in_csr_translator:av_address -> fifo_1_stage1_to_2:wrclk_control_slave_address
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_write;                                     // fifo_1_stage1_to_2_in_csr_translator:av_write -> fifo_1_stage1_to_2:wrclk_control_slave_write
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_read;                                      // fifo_1_stage1_to_2_in_csr_translator:av_read -> fifo_1_stage1_to_2:wrclk_control_slave_read
	wire   [31:0] fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_readdata;                                  // fifo_1_stage1_to_2:wrclk_control_slave_readdata -> fifo_1_stage1_to_2_in_csr_translator:av_readdata
	wire          fifo_stage1_to_4_in_translator_avalon_anti_slave_0_waitrequest;                                     // fifo_stage1_to_4:avalonmm_write_slave_waitrequest -> fifo_stage1_to_4_in_translator:av_waitrequest
	wire   [31:0] fifo_stage1_to_4_in_translator_avalon_anti_slave_0_writedata;                                       // fifo_stage1_to_4_in_translator:av_writedata -> fifo_stage1_to_4:avalonmm_write_slave_writedata
	wire          fifo_stage1_to_4_in_translator_avalon_anti_slave_0_write;                                           // fifo_stage1_to_4_in_translator:av_write -> fifo_stage1_to_4:avalonmm_write_slave_write
	wire   [31:0] fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_writedata;                                   // fifo_stage1_to_4_in_csr_translator:av_writedata -> fifo_stage1_to_4:wrclk_control_slave_writedata
	wire    [2:0] fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_address;                                     // fifo_stage1_to_4_in_csr_translator:av_address -> fifo_stage1_to_4:wrclk_control_slave_address
	wire          fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_write;                                       // fifo_stage1_to_4_in_csr_translator:av_write -> fifo_stage1_to_4:wrclk_control_slave_write
	wire          fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_read;                                        // fifo_stage1_to_4_in_csr_translator:av_read -> fifo_stage1_to_4:wrclk_control_slave_read
	wire   [31:0] fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_readdata;                                    // fifo_stage1_to_4:wrclk_control_slave_readdata -> fifo_stage1_to_4_in_csr_translator:av_readdata
	wire          fifo_stage1_to_5_in_translator_avalon_anti_slave_0_waitrequest;                                     // fifo_stage1_to_5:avalonmm_write_slave_waitrequest -> fifo_stage1_to_5_in_translator:av_waitrequest
	wire   [31:0] fifo_stage1_to_5_in_translator_avalon_anti_slave_0_writedata;                                       // fifo_stage1_to_5_in_translator:av_writedata -> fifo_stage1_to_5:avalonmm_write_slave_writedata
	wire          fifo_stage1_to_5_in_translator_avalon_anti_slave_0_write;                                           // fifo_stage1_to_5_in_translator:av_write -> fifo_stage1_to_5:avalonmm_write_slave_write
	wire   [31:0] fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_writedata;                                   // fifo_stage1_to_5_in_csr_translator:av_writedata -> fifo_stage1_to_5:wrclk_control_slave_writedata
	wire    [2:0] fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_address;                                     // fifo_stage1_to_5_in_csr_translator:av_address -> fifo_stage1_to_5:wrclk_control_slave_address
	wire          fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_write;                                       // fifo_stage1_to_5_in_csr_translator:av_write -> fifo_stage1_to_5:wrclk_control_slave_write
	wire          fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_read;                                        // fifo_stage1_to_5_in_csr_translator:av_read -> fifo_stage1_to_5:wrclk_control_slave_read
	wire   [31:0] fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_readdata;                                    // fifo_stage1_to_5:wrclk_control_slave_readdata -> fifo_stage1_to_5_in_csr_translator:av_readdata
	wire          fifo_stage1_to_6_in_translator_avalon_anti_slave_0_waitrequest;                                     // fifo_stage1_to_6:avalonmm_write_slave_waitrequest -> fifo_stage1_to_6_in_translator:av_waitrequest
	wire    [7:0] fifo_stage1_to_6_in_translator_avalon_anti_slave_0_writedata;                                       // fifo_stage1_to_6_in_translator:av_writedata -> fifo_stage1_to_6:avalonmm_write_slave_writedata
	wire          fifo_stage1_to_6_in_translator_avalon_anti_slave_0_write;                                           // fifo_stage1_to_6_in_translator:av_write -> fifo_stage1_to_6:avalonmm_write_slave_write
	wire   [31:0] fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_writedata;                                   // fifo_stage1_to_6_in_csr_translator:av_writedata -> fifo_stage1_to_6:wrclk_control_slave_writedata
	wire    [2:0] fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_address;                                     // fifo_stage1_to_6_in_csr_translator:av_address -> fifo_stage1_to_6:wrclk_control_slave_address
	wire          fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_write;                                       // fifo_stage1_to_6_in_csr_translator:av_write -> fifo_stage1_to_6:wrclk_control_slave_write
	wire          fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_read;                                        // fifo_stage1_to_6_in_csr_translator:av_read -> fifo_stage1_to_6:wrclk_control_slave_read
	wire   [31:0] fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_readdata;                                    // fifo_stage1_to_6:wrclk_control_slave_readdata -> fifo_stage1_to_6_in_csr_translator:av_readdata
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_writedata;                                             // pll_pll_slave_translator:av_writedata -> pll:writedata
	wire    [1:0] pll_pll_slave_translator_avalon_anti_slave_0_address;                                               // pll_pll_slave_translator:av_address -> pll:address
	wire          pll_pll_slave_translator_avalon_anti_slave_0_write;                                                 // pll_pll_slave_translator:av_write -> pll:write
	wire          pll_pll_slave_translator_avalon_anti_slave_0_read;                                                  // pll_pll_slave_translator:av_read -> pll:read
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_readdata;                                              // pll:readdata -> pll_pll_slave_translator:av_readdata
	wire   [31:0] instruction_mem_5_s1_translator_avalon_anti_slave_0_writedata;                                      // instruction_mem_5_s1_translator:av_writedata -> instruction_mem_5:writedata
	wire    [7:0] instruction_mem_5_s1_translator_avalon_anti_slave_0_address;                                        // instruction_mem_5_s1_translator:av_address -> instruction_mem_5:address
	wire          instruction_mem_5_s1_translator_avalon_anti_slave_0_chipselect;                                     // instruction_mem_5_s1_translator:av_chipselect -> instruction_mem_5:chipselect
	wire          instruction_mem_5_s1_translator_avalon_anti_slave_0_clken;                                          // instruction_mem_5_s1_translator:av_clken -> instruction_mem_5:clken
	wire          instruction_mem_5_s1_translator_avalon_anti_slave_0_write;                                          // instruction_mem_5_s1_translator:av_write -> instruction_mem_5:write
	wire   [31:0] instruction_mem_5_s1_translator_avalon_anti_slave_0_readdata;                                       // instruction_mem_5:readdata -> instruction_mem_5_s1_translator:av_readdata
	wire    [3:0] instruction_mem_5_s1_translator_avalon_anti_slave_0_byteenable;                                     // instruction_mem_5_s1_translator:av_byteenable -> instruction_mem_5:byteenable
	wire   [31:0] cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_5_jtag_debug_module_translator:av_writedata -> cpu_5:jtag_debug_module_writedata
	wire    [8:0] cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_5_jtag_debug_module_translator:av_address -> cpu_5:jtag_debug_module_address
	wire          cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_5_jtag_debug_module_translator:av_chipselect -> cpu_5:jtag_debug_module_select
	wire          cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_5_jtag_debug_module_translator:av_write -> cpu_5:jtag_debug_module_write
	wire   [31:0] cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_5:jtag_debug_module_readdata -> cpu_5_jtag_debug_module_translator:av_readdata
	wire          cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_5_jtag_debug_module_translator:av_begintransfer -> cpu_5:jtag_debug_module_begintransfer
	wire          cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_5_jtag_debug_module_translator:av_debugaccess -> cpu_5:jtag_debug_module_debugaccess
	wire    [3:0] cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_5_jtag_debug_module_translator:av_byteenable -> cpu_5:jtag_debug_module_byteenable
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_5:av_waitrequest -> jtag_uart_5_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_5_avalon_jtag_slave_translator:av_writedata -> jtag_uart_5:av_writedata
	wire    [0:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_5_avalon_jtag_slave_translator:av_address -> jtag_uart_5:av_address
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_5_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_5:av_chipselect
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_5_avalon_jtag_slave_translator:av_write -> jtag_uart_5:av_write_n
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_5_avalon_jtag_slave_translator:av_read -> jtag_uart_5:av_read_n
	wire   [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_5:av_readdata -> jtag_uart_5_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] timer_5_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_5_s1_translator:av_writedata -> timer_5:writedata
	wire    [2:0] timer_5_s1_translator_avalon_anti_slave_0_address;                                                  // timer_5_s1_translator:av_address -> timer_5:address
	wire          timer_5_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_5_s1_translator:av_chipselect -> timer_5:chipselect
	wire          timer_5_s1_translator_avalon_anti_slave_0_write;                                                    // timer_5_s1_translator:av_write -> timer_5:write_n
	wire   [15:0] timer_5_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_5:readdata -> timer_5_s1_translator:av_readdata
	wire          fifo_stage1_to_6_out_translator_avalon_anti_slave_0_waitrequest;                                    // fifo_stage1_to_6:avalonmm_read_slave_waitrequest -> fifo_stage1_to_6_out_translator:av_waitrequest
	wire          fifo_stage1_to_6_out_translator_avalon_anti_slave_0_read;                                           // fifo_stage1_to_6_out_translator:av_read -> fifo_stage1_to_6:avalonmm_read_slave_read
	wire    [7:0] fifo_stage1_to_6_out_translator_avalon_anti_slave_0_readdata;                                       // fifo_stage1_to_6:avalonmm_read_slave_readdata -> fifo_stage1_to_6_out_translator:av_readdata
	wire          fifo_stage5_to_6_out_translator_avalon_anti_slave_0_waitrequest;                                    // fifo_stage5_to_6:avalonmm_read_slave_waitrequest -> fifo_stage5_to_6_out_translator:av_waitrequest
	wire          fifo_stage5_to_6_out_translator_avalon_anti_slave_0_read;                                           // fifo_stage5_to_6_out_translator:av_read -> fifo_stage5_to_6:avalonmm_read_slave_read
	wire   [31:0] fifo_stage5_to_6_out_translator_avalon_anti_slave_0_readdata;                                       // fifo_stage5_to_6:avalonmm_read_slave_readdata -> fifo_stage5_to_6_out_translator:av_readdata
	wire   [31:0] fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_writedata;                                   // fifo_stage5_to_6_in_csr_translator:av_writedata -> fifo_stage5_to_6:wrclk_control_slave_writedata
	wire    [2:0] fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_address;                                     // fifo_stage5_to_6_in_csr_translator:av_address -> fifo_stage5_to_6:wrclk_control_slave_address
	wire          fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_write;                                       // fifo_stage5_to_6_in_csr_translator:av_write -> fifo_stage5_to_6:wrclk_control_slave_write
	wire          fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_read;                                        // fifo_stage5_to_6_in_csr_translator:av_read -> fifo_stage5_to_6:wrclk_control_slave_read
	wire   [31:0] fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_readdata;                                    // fifo_stage5_to_6:wrclk_control_slave_readdata -> fifo_stage5_to_6_in_csr_translator:av_readdata
	wire   [31:0] instruction_mem_1_s1_translator_avalon_anti_slave_0_writedata;                                      // instruction_mem_1_s1_translator:av_writedata -> instruction_mem_1:writedata
	wire    [7:0] instruction_mem_1_s1_translator_avalon_anti_slave_0_address;                                        // instruction_mem_1_s1_translator:av_address -> instruction_mem_1:address
	wire          instruction_mem_1_s1_translator_avalon_anti_slave_0_chipselect;                                     // instruction_mem_1_s1_translator:av_chipselect -> instruction_mem_1:chipselect
	wire          instruction_mem_1_s1_translator_avalon_anti_slave_0_clken;                                          // instruction_mem_1_s1_translator:av_clken -> instruction_mem_1:clken
	wire          instruction_mem_1_s1_translator_avalon_anti_slave_0_write;                                          // instruction_mem_1_s1_translator:av_write -> instruction_mem_1:write
	wire   [31:0] instruction_mem_1_s1_translator_avalon_anti_slave_0_readdata;                                       // instruction_mem_1:readdata -> instruction_mem_1_s1_translator:av_readdata
	wire    [3:0] instruction_mem_1_s1_translator_avalon_anti_slave_0_byteenable;                                     // instruction_mem_1_s1_translator:av_byteenable -> instruction_mem_1:byteenable
	wire   [31:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_1_jtag_debug_module_translator:av_writedata -> cpu_1:jtag_debug_module_writedata
	wire    [8:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_1_jtag_debug_module_translator:av_address -> cpu_1:jtag_debug_module_address
	wire          cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_1_jtag_debug_module_translator:av_chipselect -> cpu_1:jtag_debug_module_select
	wire          cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_1_jtag_debug_module_translator:av_write -> cpu_1:jtag_debug_module_write
	wire   [31:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_1:jtag_debug_module_readdata -> cpu_1_jtag_debug_module_translator:av_readdata
	wire          cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_1_jtag_debug_module_translator:av_begintransfer -> cpu_1:jtag_debug_module_begintransfer
	wire          cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_1_jtag_debug_module_translator:av_debugaccess -> cpu_1:jtag_debug_module_debugaccess
	wire    [3:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_1_jtag_debug_module_translator:av_byteenable -> cpu_1:jtag_debug_module_byteenable
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_1:av_waitrequest -> jtag_uart_1_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_1_avalon_jtag_slave_translator:av_writedata -> jtag_uart_1:av_writedata
	wire    [0:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_1_avalon_jtag_slave_translator:av_address -> jtag_uart_1:av_address
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_1_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_1:av_chipselect
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_1_avalon_jtag_slave_translator:av_write -> jtag_uart_1:av_write_n
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_1_avalon_jtag_slave_translator:av_read -> jtag_uart_1:av_read_n
	wire   [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_1:av_readdata -> jtag_uart_1_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] timer_1_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_1_s1_translator:av_writedata -> timer_1:writedata
	wire    [2:0] timer_1_s1_translator_avalon_anti_slave_0_address;                                                  // timer_1_s1_translator:av_address -> timer_1:address
	wire          timer_1_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	wire          timer_1_s1_translator_avalon_anti_slave_0_write;                                                    // timer_1_s1_translator:av_write -> timer_1:write_n
	wire   [15:0] timer_1_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_1:readdata -> timer_1_s1_translator:av_readdata
	wire          fifo_0_stage1_to_2_out_translator_avalon_anti_slave_0_waitrequest;                                  // fifo_0_stage1_to_2:avalonmm_read_slave_waitrequest -> fifo_0_stage1_to_2_out_translator:av_waitrequest
	wire          fifo_0_stage1_to_2_out_translator_avalon_anti_slave_0_read;                                         // fifo_0_stage1_to_2_out_translator:av_read -> fifo_0_stage1_to_2:avalonmm_read_slave_read
	wire   [31:0] fifo_0_stage1_to_2_out_translator_avalon_anti_slave_0_readdata;                                     // fifo_0_stage1_to_2:avalonmm_read_slave_readdata -> fifo_0_stage1_to_2_out_translator:av_readdata
	wire          fifo_1_stage1_to_2_out_translator_avalon_anti_slave_0_waitrequest;                                  // fifo_1_stage1_to_2:avalonmm_read_slave_waitrequest -> fifo_1_stage1_to_2_out_translator:av_waitrequest
	wire          fifo_1_stage1_to_2_out_translator_avalon_anti_slave_0_read;                                         // fifo_1_stage1_to_2_out_translator:av_read -> fifo_1_stage1_to_2:avalonmm_read_slave_read
	wire   [31:0] fifo_1_stage1_to_2_out_translator_avalon_anti_slave_0_readdata;                                     // fifo_1_stage1_to_2:avalonmm_read_slave_readdata -> fifo_1_stage1_to_2_out_translator:av_readdata
	wire          fifo_2_stage1_to_2_out_translator_avalon_anti_slave_0_waitrequest;                                  // fifo_2_stage1_to_2:avalonmm_read_slave_waitrequest -> fifo_2_stage1_to_2_out_translator:av_waitrequest
	wire          fifo_2_stage1_to_2_out_translator_avalon_anti_slave_0_read;                                         // fifo_2_stage1_to_2_out_translator:av_read -> fifo_2_stage1_to_2:avalonmm_read_slave_read
	wire   [31:0] fifo_2_stage1_to_2_out_translator_avalon_anti_slave_0_readdata;                                     // fifo_2_stage1_to_2:avalonmm_read_slave_readdata -> fifo_2_stage1_to_2_out_translator:av_readdata
	wire          fifo_stage2_to_3_in_translator_avalon_anti_slave_0_waitrequest;                                     // fifo_stage2_to_3:avalonmm_write_slave_waitrequest -> fifo_stage2_to_3_in_translator:av_waitrequest
	wire   [31:0] fifo_stage2_to_3_in_translator_avalon_anti_slave_0_writedata;                                       // fifo_stage2_to_3_in_translator:av_writedata -> fifo_stage2_to_3:avalonmm_write_slave_writedata
	wire          fifo_stage2_to_3_in_translator_avalon_anti_slave_0_write;                                           // fifo_stage2_to_3_in_translator:av_write -> fifo_stage2_to_3:avalonmm_write_slave_write
	wire   [31:0] fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_writedata;                                   // fifo_stage2_to_3_in_csr_translator:av_writedata -> fifo_stage2_to_3:wrclk_control_slave_writedata
	wire    [2:0] fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_address;                                     // fifo_stage2_to_3_in_csr_translator:av_address -> fifo_stage2_to_3:wrclk_control_slave_address
	wire          fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_write;                                       // fifo_stage2_to_3_in_csr_translator:av_write -> fifo_stage2_to_3:wrclk_control_slave_write
	wire          fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_read;                                        // fifo_stage2_to_3_in_csr_translator:av_read -> fifo_stage2_to_3:wrclk_control_slave_read
	wire   [31:0] fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_readdata;                                    // fifo_stage2_to_3:wrclk_control_slave_readdata -> fifo_stage2_to_3_in_csr_translator:av_readdata
	wire   [31:0] instruction_mem_2_s1_translator_avalon_anti_slave_0_writedata;                                      // instruction_mem_2_s1_translator:av_writedata -> instruction_mem_2:writedata
	wire    [7:0] instruction_mem_2_s1_translator_avalon_anti_slave_0_address;                                        // instruction_mem_2_s1_translator:av_address -> instruction_mem_2:address
	wire          instruction_mem_2_s1_translator_avalon_anti_slave_0_chipselect;                                     // instruction_mem_2_s1_translator:av_chipselect -> instruction_mem_2:chipselect
	wire          instruction_mem_2_s1_translator_avalon_anti_slave_0_clken;                                          // instruction_mem_2_s1_translator:av_clken -> instruction_mem_2:clken
	wire          instruction_mem_2_s1_translator_avalon_anti_slave_0_write;                                          // instruction_mem_2_s1_translator:av_write -> instruction_mem_2:write
	wire   [31:0] instruction_mem_2_s1_translator_avalon_anti_slave_0_readdata;                                       // instruction_mem_2:readdata -> instruction_mem_2_s1_translator:av_readdata
	wire    [3:0] instruction_mem_2_s1_translator_avalon_anti_slave_0_byteenable;                                     // instruction_mem_2_s1_translator:av_byteenable -> instruction_mem_2:byteenable
	wire   [31:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_2_jtag_debug_module_translator:av_writedata -> cpu_2:jtag_debug_module_writedata
	wire    [8:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_2_jtag_debug_module_translator:av_address -> cpu_2:jtag_debug_module_address
	wire          cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_2_jtag_debug_module_translator:av_chipselect -> cpu_2:jtag_debug_module_select
	wire          cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_2_jtag_debug_module_translator:av_write -> cpu_2:jtag_debug_module_write
	wire   [31:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_2:jtag_debug_module_readdata -> cpu_2_jtag_debug_module_translator:av_readdata
	wire          cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_2_jtag_debug_module_translator:av_begintransfer -> cpu_2:jtag_debug_module_begintransfer
	wire          cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_2_jtag_debug_module_translator:av_debugaccess -> cpu_2:jtag_debug_module_debugaccess
	wire    [3:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_2_jtag_debug_module_translator:av_byteenable -> cpu_2:jtag_debug_module_byteenable
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_2:av_waitrequest -> jtag_uart_2_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_2_avalon_jtag_slave_translator:av_writedata -> jtag_uart_2:av_writedata
	wire    [0:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_2_avalon_jtag_slave_translator:av_address -> jtag_uart_2:av_address
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_2_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_2:av_chipselect
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_2_avalon_jtag_slave_translator:av_write -> jtag_uart_2:av_write_n
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_2_avalon_jtag_slave_translator:av_read -> jtag_uart_2:av_read_n
	wire   [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_2:av_readdata -> jtag_uart_2_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] timer_2_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_2_s1_translator:av_writedata -> timer_2:writedata
	wire    [2:0] timer_2_s1_translator_avalon_anti_slave_0_address;                                                  // timer_2_s1_translator:av_address -> timer_2:address
	wire          timer_2_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_2_s1_translator:av_chipselect -> timer_2:chipselect
	wire          timer_2_s1_translator_avalon_anti_slave_0_write;                                                    // timer_2_s1_translator:av_write -> timer_2:write_n
	wire   [15:0] timer_2_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_2:readdata -> timer_2_s1_translator:av_readdata
	wire          fifo_stage2_to_3_out_translator_avalon_anti_slave_0_waitrequest;                                    // fifo_stage2_to_3:avalonmm_read_slave_waitrequest -> fifo_stage2_to_3_out_translator:av_waitrequest
	wire          fifo_stage2_to_3_out_translator_avalon_anti_slave_0_read;                                           // fifo_stage2_to_3_out_translator:av_read -> fifo_stage2_to_3:avalonmm_read_slave_read
	wire   [31:0] fifo_stage2_to_3_out_translator_avalon_anti_slave_0_readdata;                                       // fifo_stage2_to_3:avalonmm_read_slave_readdata -> fifo_stage2_to_3_out_translator:av_readdata
	wire          fifo_stage3_to_4_in_translator_avalon_anti_slave_0_waitrequest;                                     // fifo_stage3_to_4:avalonmm_write_slave_waitrequest -> fifo_stage3_to_4_in_translator:av_waitrequest
	wire   [31:0] fifo_stage3_to_4_in_translator_avalon_anti_slave_0_writedata;                                       // fifo_stage3_to_4_in_translator:av_writedata -> fifo_stage3_to_4:avalonmm_write_slave_writedata
	wire          fifo_stage3_to_4_in_translator_avalon_anti_slave_0_write;                                           // fifo_stage3_to_4_in_translator:av_write -> fifo_stage3_to_4:avalonmm_write_slave_write
	wire   [31:0] fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_writedata;                                   // fifo_stage3_to_4_in_csr_translator:av_writedata -> fifo_stage3_to_4:wrclk_control_slave_writedata
	wire    [2:0] fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_address;                                     // fifo_stage3_to_4_in_csr_translator:av_address -> fifo_stage3_to_4:wrclk_control_slave_address
	wire          fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_write;                                       // fifo_stage3_to_4_in_csr_translator:av_write -> fifo_stage3_to_4:wrclk_control_slave_write
	wire          fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_read;                                        // fifo_stage3_to_4_in_csr_translator:av_read -> fifo_stage3_to_4:wrclk_control_slave_read
	wire   [31:0] fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_readdata;                                    // fifo_stage3_to_4:wrclk_control_slave_readdata -> fifo_stage3_to_4_in_csr_translator:av_readdata
	wire   [31:0] instruction_mem_3_s1_translator_avalon_anti_slave_0_writedata;                                      // instruction_mem_3_s1_translator:av_writedata -> instruction_mem_3:writedata
	wire    [7:0] instruction_mem_3_s1_translator_avalon_anti_slave_0_address;                                        // instruction_mem_3_s1_translator:av_address -> instruction_mem_3:address
	wire          instruction_mem_3_s1_translator_avalon_anti_slave_0_chipselect;                                     // instruction_mem_3_s1_translator:av_chipselect -> instruction_mem_3:chipselect
	wire          instruction_mem_3_s1_translator_avalon_anti_slave_0_clken;                                          // instruction_mem_3_s1_translator:av_clken -> instruction_mem_3:clken
	wire          instruction_mem_3_s1_translator_avalon_anti_slave_0_write;                                          // instruction_mem_3_s1_translator:av_write -> instruction_mem_3:write
	wire   [31:0] instruction_mem_3_s1_translator_avalon_anti_slave_0_readdata;                                       // instruction_mem_3:readdata -> instruction_mem_3_s1_translator:av_readdata
	wire    [3:0] instruction_mem_3_s1_translator_avalon_anti_slave_0_byteenable;                                     // instruction_mem_3_s1_translator:av_byteenable -> instruction_mem_3:byteenable
	wire   [31:0] cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_3_jtag_debug_module_translator:av_writedata -> cpu_3:jtag_debug_module_writedata
	wire    [8:0] cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_3_jtag_debug_module_translator:av_address -> cpu_3:jtag_debug_module_address
	wire          cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_3_jtag_debug_module_translator:av_chipselect -> cpu_3:jtag_debug_module_select
	wire          cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_3_jtag_debug_module_translator:av_write -> cpu_3:jtag_debug_module_write
	wire   [31:0] cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_3:jtag_debug_module_readdata -> cpu_3_jtag_debug_module_translator:av_readdata
	wire          cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_3_jtag_debug_module_translator:av_begintransfer -> cpu_3:jtag_debug_module_begintransfer
	wire          cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_3_jtag_debug_module_translator:av_debugaccess -> cpu_3:jtag_debug_module_debugaccess
	wire    [3:0] cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_3_jtag_debug_module_translator:av_byteenable -> cpu_3:jtag_debug_module_byteenable
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_3:av_waitrequest -> jtag_uart_3_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_3_avalon_jtag_slave_translator:av_writedata -> jtag_uart_3:av_writedata
	wire    [0:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_3_avalon_jtag_slave_translator:av_address -> jtag_uart_3:av_address
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_3_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_3:av_chipselect
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_3_avalon_jtag_slave_translator:av_write -> jtag_uart_3:av_write_n
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_3_avalon_jtag_slave_translator:av_read -> jtag_uart_3:av_read_n
	wire   [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_3:av_readdata -> jtag_uart_3_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] timer_3_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_3_s1_translator:av_writedata -> timer_3:writedata
	wire    [2:0] timer_3_s1_translator_avalon_anti_slave_0_address;                                                  // timer_3_s1_translator:av_address -> timer_3:address
	wire          timer_3_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_3_s1_translator:av_chipselect -> timer_3:chipselect
	wire          timer_3_s1_translator_avalon_anti_slave_0_write;                                                    // timer_3_s1_translator:av_write -> timer_3:write_n
	wire   [15:0] timer_3_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_3:readdata -> timer_3_s1_translator:av_readdata
	wire          fifo_stage1_to_4_out_translator_avalon_anti_slave_0_waitrequest;                                    // fifo_stage1_to_4:avalonmm_read_slave_waitrequest -> fifo_stage1_to_4_out_translator:av_waitrequest
	wire          fifo_stage1_to_4_out_translator_avalon_anti_slave_0_read;                                           // fifo_stage1_to_4_out_translator:av_read -> fifo_stage1_to_4:avalonmm_read_slave_read
	wire   [31:0] fifo_stage1_to_4_out_translator_avalon_anti_slave_0_readdata;                                       // fifo_stage1_to_4:avalonmm_read_slave_readdata -> fifo_stage1_to_4_out_translator:av_readdata
	wire          fifo_stage3_to_4_out_translator_avalon_anti_slave_0_waitrequest;                                    // fifo_stage3_to_4:avalonmm_read_slave_waitrequest -> fifo_stage3_to_4_out_translator:av_waitrequest
	wire          fifo_stage3_to_4_out_translator_avalon_anti_slave_0_read;                                           // fifo_stage3_to_4_out_translator:av_read -> fifo_stage3_to_4:avalonmm_read_slave_read
	wire   [31:0] fifo_stage3_to_4_out_translator_avalon_anti_slave_0_readdata;                                       // fifo_stage3_to_4:avalonmm_read_slave_readdata -> fifo_stage3_to_4_out_translator:av_readdata
	wire          fifo_stage4_to_5_in_translator_avalon_anti_slave_0_waitrequest;                                     // fifo_stage4_to_5:avalonmm_write_slave_waitrequest -> fifo_stage4_to_5_in_translator:av_waitrequest
	wire   [31:0] fifo_stage4_to_5_in_translator_avalon_anti_slave_0_writedata;                                       // fifo_stage4_to_5_in_translator:av_writedata -> fifo_stage4_to_5:avalonmm_write_slave_writedata
	wire          fifo_stage4_to_5_in_translator_avalon_anti_slave_0_write;                                           // fifo_stage4_to_5_in_translator:av_write -> fifo_stage4_to_5:avalonmm_write_slave_write
	wire   [31:0] fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_writedata;                                   // fifo_stage4_to_5_in_csr_translator:av_writedata -> fifo_stage4_to_5:wrclk_control_slave_writedata
	wire    [2:0] fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_address;                                     // fifo_stage4_to_5_in_csr_translator:av_address -> fifo_stage4_to_5:wrclk_control_slave_address
	wire          fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_write;                                       // fifo_stage4_to_5_in_csr_translator:av_write -> fifo_stage4_to_5:wrclk_control_slave_write
	wire          fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_read;                                        // fifo_stage4_to_5_in_csr_translator:av_read -> fifo_stage4_to_5:wrclk_control_slave_read
	wire   [31:0] fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_readdata;                                    // fifo_stage4_to_5:wrclk_control_slave_readdata -> fifo_stage4_to_5_in_csr_translator:av_readdata
	wire   [31:0] instruction_mem_4_s1_translator_avalon_anti_slave_0_writedata;                                      // instruction_mem_4_s1_translator:av_writedata -> instruction_mem_4:writedata
	wire    [7:0] instruction_mem_4_s1_translator_avalon_anti_slave_0_address;                                        // instruction_mem_4_s1_translator:av_address -> instruction_mem_4:address
	wire          instruction_mem_4_s1_translator_avalon_anti_slave_0_chipselect;                                     // instruction_mem_4_s1_translator:av_chipselect -> instruction_mem_4:chipselect
	wire          instruction_mem_4_s1_translator_avalon_anti_slave_0_clken;                                          // instruction_mem_4_s1_translator:av_clken -> instruction_mem_4:clken
	wire          instruction_mem_4_s1_translator_avalon_anti_slave_0_write;                                          // instruction_mem_4_s1_translator:av_write -> instruction_mem_4:write
	wire   [31:0] instruction_mem_4_s1_translator_avalon_anti_slave_0_readdata;                                       // instruction_mem_4:readdata -> instruction_mem_4_s1_translator:av_readdata
	wire    [3:0] instruction_mem_4_s1_translator_avalon_anti_slave_0_byteenable;                                     // instruction_mem_4_s1_translator:av_byteenable -> instruction_mem_4:byteenable
	wire   [31:0] cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_4_jtag_debug_module_translator:av_writedata -> cpu_4:jtag_debug_module_writedata
	wire    [8:0] cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_4_jtag_debug_module_translator:av_address -> cpu_4:jtag_debug_module_address
	wire          cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_4_jtag_debug_module_translator:av_chipselect -> cpu_4:jtag_debug_module_select
	wire          cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_4_jtag_debug_module_translator:av_write -> cpu_4:jtag_debug_module_write
	wire   [31:0] cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_4:jtag_debug_module_readdata -> cpu_4_jtag_debug_module_translator:av_readdata
	wire          cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_4_jtag_debug_module_translator:av_begintransfer -> cpu_4:jtag_debug_module_begintransfer
	wire          cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_4_jtag_debug_module_translator:av_debugaccess -> cpu_4:jtag_debug_module_debugaccess
	wire    [3:0] cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_4_jtag_debug_module_translator:av_byteenable -> cpu_4:jtag_debug_module_byteenable
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_4:av_waitrequest -> jtag_uart_4_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_4_avalon_jtag_slave_translator:av_writedata -> jtag_uart_4:av_writedata
	wire    [0:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_4_avalon_jtag_slave_translator:av_address -> jtag_uart_4:av_address
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_4_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_4:av_chipselect
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_4_avalon_jtag_slave_translator:av_write -> jtag_uart_4:av_write_n
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_4_avalon_jtag_slave_translator:av_read -> jtag_uart_4:av_read_n
	wire   [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_4:av_readdata -> jtag_uart_4_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] timer_4_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_4_s1_translator:av_writedata -> timer_4:writedata
	wire    [2:0] timer_4_s1_translator_avalon_anti_slave_0_address;                                                  // timer_4_s1_translator:av_address -> timer_4:address
	wire          timer_4_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_4_s1_translator:av_chipselect -> timer_4:chipselect
	wire          timer_4_s1_translator_avalon_anti_slave_0_write;                                                    // timer_4_s1_translator:av_write -> timer_4:write_n
	wire   [15:0] timer_4_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_4:readdata -> timer_4_s1_translator:av_readdata
	wire          fifo_stage1_to_5_out_translator_avalon_anti_slave_0_waitrequest;                                    // fifo_stage1_to_5:avalonmm_read_slave_waitrequest -> fifo_stage1_to_5_out_translator:av_waitrequest
	wire          fifo_stage1_to_5_out_translator_avalon_anti_slave_0_read;                                           // fifo_stage1_to_5_out_translator:av_read -> fifo_stage1_to_5:avalonmm_read_slave_read
	wire   [31:0] fifo_stage1_to_5_out_translator_avalon_anti_slave_0_readdata;                                       // fifo_stage1_to_5:avalonmm_read_slave_readdata -> fifo_stage1_to_5_out_translator:av_readdata
	wire          fifo_stage4_to_5_out_translator_avalon_anti_slave_0_waitrequest;                                    // fifo_stage4_to_5:avalonmm_read_slave_waitrequest -> fifo_stage4_to_5_out_translator:av_waitrequest
	wire          fifo_stage4_to_5_out_translator_avalon_anti_slave_0_read;                                           // fifo_stage4_to_5_out_translator:av_read -> fifo_stage4_to_5:avalonmm_read_slave_read
	wire   [31:0] fifo_stage4_to_5_out_translator_avalon_anti_slave_0_readdata;                                       // fifo_stage4_to_5:avalonmm_read_slave_readdata -> fifo_stage4_to_5_out_translator:av_readdata
	wire          fifo_stage5_to_6_in_translator_avalon_anti_slave_0_waitrequest;                                     // fifo_stage5_to_6:avalonmm_write_slave_waitrequest -> fifo_stage5_to_6_in_translator:av_waitrequest
	wire   [31:0] fifo_stage5_to_6_in_translator_avalon_anti_slave_0_writedata;                                       // fifo_stage5_to_6_in_translator:av_writedata -> fifo_stage5_to_6:avalonmm_write_slave_writedata
	wire          fifo_stage5_to_6_in_translator_avalon_anti_slave_0_write;                                           // fifo_stage5_to_6_in_translator:av_write -> fifo_stage5_to_6:avalonmm_write_slave_write
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_0_instruction_master_translator:uav_burstcount -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_0_instruction_master_translator:uav_writedata -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_0_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_0_instruction_master_translator:uav_address -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_0_instruction_master_translator:uav_lock -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_0_instruction_master_translator:uav_write -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_0_instruction_master_translator:uav_read -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_instruction_master_translator:uav_readdata
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_0_instruction_master_translator:uav_debugaccess -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_0_instruction_master_translator:uav_byteenable -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_instruction_master_translator:uav_readdatavalid
	wire          cpu_0_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_0_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_0_data_master_translator:uav_burstcount -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_0_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_0_data_master_translator:uav_writedata -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_0_data_master_translator_avalon_universal_master_0_address;                                     // cpu_0_data_master_translator:uav_address -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_0_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_0_data_master_translator:uav_lock -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_0_data_master_translator_avalon_universal_master_0_write;                                       // cpu_0_data_master_translator:uav_write -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_0_data_master_translator_avalon_universal_master_0_read;                                        // cpu_0_data_master_translator:uav_read -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_0_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_data_master_translator:uav_readdata
	wire          cpu_0_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_0_data_master_translator:uav_debugaccess -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_0_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_0_data_master_translator:uav_byteenable -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_data_master_translator:uav_readdatavalid
	wire          cpu_5_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_5_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_5_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_5_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_5_data_master_translator:uav_burstcount -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_5_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_5_data_master_translator:uav_writedata -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_5_data_master_translator_avalon_universal_master_0_address;                                     // cpu_5_data_master_translator:uav_address -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_5_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_5_data_master_translator:uav_lock -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_5_data_master_translator_avalon_universal_master_0_write;                                       // cpu_5_data_master_translator:uav_write -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_5_data_master_translator_avalon_universal_master_0_read;                                        // cpu_5_data_master_translator:uav_read -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_5_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_5_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_5_data_master_translator:uav_readdata
	wire          cpu_5_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_5_data_master_translator:uav_debugaccess -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_5_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_5_data_master_translator:uav_byteenable -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_5_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_5_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_5_data_master_translator:uav_readdatavalid
	wire          cpu_4_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_4_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_4_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_4_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_4_data_master_translator:uav_burstcount -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_4_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_4_data_master_translator:uav_writedata -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_4_data_master_translator_avalon_universal_master_0_address;                                     // cpu_4_data_master_translator:uav_address -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_4_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_4_data_master_translator:uav_lock -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_4_data_master_translator_avalon_universal_master_0_write;                                       // cpu_4_data_master_translator:uav_write -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_4_data_master_translator_avalon_universal_master_0_read;                                        // cpu_4_data_master_translator:uav_read -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_4_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_4_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_4_data_master_translator:uav_readdata
	wire          cpu_4_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_4_data_master_translator:uav_debugaccess -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_4_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_4_data_master_translator:uav_byteenable -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_4_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_4_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_4_data_master_translator:uav_readdatavalid
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_4_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_4_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_4_instruction_master_translator:uav_burstcount -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_4_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_4_instruction_master_translator:uav_writedata -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_4_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_4_instruction_master_translator:uav_address -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_4_instruction_master_translator:uav_lock -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_4_instruction_master_translator:uav_write -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_4_instruction_master_translator:uav_read -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_4_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_4_instruction_master_translator:uav_readdata
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_4_instruction_master_translator:uav_debugaccess -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_4_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_4_instruction_master_translator:uav_byteenable -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_4_instruction_master_translator:uav_readdatavalid
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_1_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_1_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_1_instruction_master_translator:uav_burstcount -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_1_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_1_instruction_master_translator:uav_writedata -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_1_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_1_instruction_master_translator:uav_address -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_1_instruction_master_translator:uav_lock -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_1_instruction_master_translator:uav_write -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_1_instruction_master_translator:uav_read -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_1_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_1_instruction_master_translator:uav_readdata
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_1_instruction_master_translator:uav_debugaccess -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_1_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_1_instruction_master_translator:uav_byteenable -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_1_instruction_master_translator:uav_readdatavalid
	wire          cpu_1_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_1_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_1_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_1_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_1_data_master_translator:uav_burstcount -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_1_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_1_data_master_translator:uav_writedata -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_1_data_master_translator_avalon_universal_master_0_address;                                     // cpu_1_data_master_translator:uav_address -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_1_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_1_data_master_translator:uav_lock -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_1_data_master_translator_avalon_universal_master_0_write;                                       // cpu_1_data_master_translator:uav_write -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_1_data_master_translator_avalon_universal_master_0_read;                                        // cpu_1_data_master_translator:uav_read -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_1_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_1_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_1_data_master_translator:uav_readdata
	wire          cpu_1_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_1_data_master_translator:uav_debugaccess -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_1_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_1_data_master_translator:uav_byteenable -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_1_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_1_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_1_data_master_translator:uav_readdatavalid
	wire          cpu_2_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_2_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_2_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_2_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_2_data_master_translator:uav_burstcount -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_2_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_2_data_master_translator:uav_writedata -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_2_data_master_translator_avalon_universal_master_0_address;                                     // cpu_2_data_master_translator:uav_address -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_2_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_2_data_master_translator:uav_lock -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_2_data_master_translator_avalon_universal_master_0_write;                                       // cpu_2_data_master_translator:uav_write -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_2_data_master_translator_avalon_universal_master_0_read;                                        // cpu_2_data_master_translator:uav_read -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_2_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_2_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_2_data_master_translator:uav_readdata
	wire          cpu_2_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_2_data_master_translator:uav_debugaccess -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_2_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_2_data_master_translator:uav_byteenable -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_2_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_2_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_2_data_master_translator:uav_readdatavalid
	wire          cpu_3_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_3_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_3_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_3_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_3_data_master_translator:uav_burstcount -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_3_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_3_data_master_translator:uav_writedata -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_3_data_master_translator_avalon_universal_master_0_address;                                     // cpu_3_data_master_translator:uav_address -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_3_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_3_data_master_translator:uav_lock -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_3_data_master_translator_avalon_universal_master_0_write;                                       // cpu_3_data_master_translator:uav_write -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_3_data_master_translator_avalon_universal_master_0_read;                                        // cpu_3_data_master_translator:uav_read -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_3_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_3_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_3_data_master_translator:uav_readdata
	wire          cpu_3_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_3_data_master_translator:uav_debugaccess -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_3_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_3_data_master_translator:uav_byteenable -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_3_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_3_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_3_data_master_translator:uav_readdatavalid
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_3_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_3_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_3_instruction_master_translator:uav_burstcount -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_3_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_3_instruction_master_translator:uav_writedata -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_3_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_3_instruction_master_translator:uav_address -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_3_instruction_master_translator:uav_lock -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_3_instruction_master_translator:uav_write -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_3_instruction_master_translator:uav_read -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_3_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_3_instruction_master_translator:uav_readdata
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_3_instruction_master_translator:uav_debugaccess -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_3_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_3_instruction_master_translator:uav_byteenable -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_3_instruction_master_translator:uav_readdatavalid
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_2_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_2_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_2_instruction_master_translator:uav_burstcount -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_2_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_2_instruction_master_translator:uav_writedata -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_2_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_2_instruction_master_translator:uav_address -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_2_instruction_master_translator:uav_lock -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_2_instruction_master_translator:uav_write -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_2_instruction_master_translator:uav_read -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_2_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_2_instruction_master_translator:uav_readdata
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_2_instruction_master_translator:uav_debugaccess -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_2_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_2_instruction_master_translator:uav_byteenable -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_2_instruction_master_translator:uav_readdatavalid
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_5_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_5_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_5_instruction_master_translator:uav_burstcount -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_5_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_5_instruction_master_translator:uav_writedata -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_5_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_5_instruction_master_translator:uav_address -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_5_instruction_master_translator:uav_lock -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_5_instruction_master_translator:uav_write -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_5_instruction_master_translator:uav_read -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_5_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_5_instruction_master_translator:uav_readdata
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_5_instruction_master_translator:uav_debugaccess -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_5_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_5_instruction_master_translator:uav_byteenable -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_5_instruction_master_translator:uav_readdatavalid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_0_jtag_debug_module_translator:uav_waitrequest -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_0_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_0_jtag_debug_module_translator:uav_writedata
	wire   [27:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_0_jtag_debug_module_translator:uav_address
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_0_jtag_debug_module_translator:uav_write
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_0_jtag_debug_module_translator:uav_lock
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_0_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_0_jtag_debug_module_translator:uav_readdata -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_0_jtag_debug_module_translator:uav_readdatavalid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_0_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_0_jtag_debug_module_translator:uav_byteenable
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // sdram_controller_s1_translator:uav_waitrequest -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_controller_s1_translator:uav_burstcount
	wire   [31:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_controller_s1_translator:uav_writedata
	wire   [27:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_controller_s1_translator:uav_address
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_controller_s1_translator:uav_write
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_controller_s1_translator:uav_lock
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_controller_s1_translator:uav_read
	wire   [31:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // sdram_controller_s1_translator:uav_readdata -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // sdram_controller_s1_translator:uav_readdatavalid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_controller_s1_translator:uav_debugaccess
	wire    [3:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_controller_s1_translator:uav_byteenable
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire   [27:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire    [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [27:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // fifo_0_stage1_to_2_in_translator:uav_waitrequest -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_stage1_to_2_in_translator:uav_burstcount
	wire   [31:0] fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata;                       // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_stage1_to_2_in_translator:uav_writedata
	wire   [27:0] fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address;                         // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_stage1_to_2_in_translator:uav_address
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write;                           // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_stage1_to_2_in_translator:uav_write
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock;                            // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_stage1_to_2_in_translator:uav_lock
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read;                            // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_stage1_to_2_in_translator:uav_read
	wire   [31:0] fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata;                        // fifo_0_stage1_to_2_in_translator:uav_readdata -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // fifo_0_stage1_to_2_in_translator:uav_readdatavalid -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_stage1_to_2_in_translator:uav_debugaccess
	wire    [3:0] fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_stage1_to_2_in_translator:uav_byteenable
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data;                     // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // fifo_0_stage1_to_2_in_csr_translator:uav_waitrequest -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_stage1_to_2_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                   // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_stage1_to_2_in_csr_translator:uav_writedata
	wire   [27:0] fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                     // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_stage1_to_2_in_csr_translator:uav_address
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                       // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_stage1_to_2_in_csr_translator:uav_write
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                        // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_stage1_to_2_in_csr_translator:uav_lock
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                        // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_stage1_to_2_in_csr_translator:uav_read
	wire   [31:0] fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                    // fifo_0_stage1_to_2_in_csr_translator:uav_readdata -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // fifo_0_stage1_to_2_in_csr_translator:uav_readdatavalid -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_stage1_to_2_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_stage1_to_2_in_csr_translator:uav_byteenable
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                 // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // fifo_1_stage1_to_2_in_translator:uav_waitrequest -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_stage1_to_2_in_translator:uav_burstcount
	wire   [31:0] fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata;                       // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_stage1_to_2_in_translator:uav_writedata
	wire   [27:0] fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address;                         // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_stage1_to_2_in_translator:uav_address
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write;                           // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_stage1_to_2_in_translator:uav_write
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock;                            // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_stage1_to_2_in_translator:uav_lock
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read;                            // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_stage1_to_2_in_translator:uav_read
	wire   [31:0] fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata;                        // fifo_1_stage1_to_2_in_translator:uav_readdata -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // fifo_1_stage1_to_2_in_translator:uav_readdatavalid -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_stage1_to_2_in_translator:uav_debugaccess
	wire    [3:0] fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_stage1_to_2_in_translator:uav_byteenable
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data;                     // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // fifo_2_stage1_to_2_in_translator:uav_waitrequest -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_stage1_to_2_in_translator:uav_burstcount
	wire   [31:0] fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata;                       // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_stage1_to_2_in_translator:uav_writedata
	wire   [27:0] fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address;                         // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_stage1_to_2_in_translator:uav_address
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write;                           // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_stage1_to_2_in_translator:uav_write
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock;                            // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_stage1_to_2_in_translator:uav_lock
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read;                            // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_stage1_to_2_in_translator:uav_read
	wire   [31:0] fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata;                        // fifo_2_stage1_to_2_in_translator:uav_readdata -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // fifo_2_stage1_to_2_in_translator:uav_readdatavalid -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_stage1_to_2_in_translator:uav_debugaccess
	wire    [3:0] fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_stage1_to_2_in_translator:uav_byteenable
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data;                     // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // fifo_2_stage1_to_2_in_csr_translator:uav_waitrequest -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_stage1_to_2_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                   // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_stage1_to_2_in_csr_translator:uav_writedata
	wire   [27:0] fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                     // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_stage1_to_2_in_csr_translator:uav_address
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                       // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_stage1_to_2_in_csr_translator:uav_write
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                        // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_stage1_to_2_in_csr_translator:uav_lock
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                        // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_stage1_to_2_in_csr_translator:uav_read
	wire   [31:0] fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                    // fifo_2_stage1_to_2_in_csr_translator:uav_readdata -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // fifo_2_stage1_to_2_in_csr_translator:uav_readdatavalid -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_stage1_to_2_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_stage1_to_2_in_csr_translator:uav_byteenable
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                 // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // fifo_1_stage1_to_2_in_csr_translator:uav_waitrequest -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_stage1_to_2_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                   // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_stage1_to_2_in_csr_translator:uav_writedata
	wire   [27:0] fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                     // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_stage1_to_2_in_csr_translator:uav_address
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                       // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_stage1_to_2_in_csr_translator:uav_write
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                        // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_stage1_to_2_in_csr_translator:uav_lock
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                        // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_stage1_to_2_in_csr_translator:uav_read
	wire   [31:0] fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                    // fifo_1_stage1_to_2_in_csr_translator:uav_readdata -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // fifo_1_stage1_to_2_in_csr_translator:uav_readdatavalid -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_stage1_to_2_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_stage1_to_2_in_csr_translator:uav_byteenable
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                 // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // fifo_stage1_to_4_in_translator:uav_waitrequest -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage1_to_4_in_translator:uav_burstcount
	wire   [31:0] fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_writedata;                         // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage1_to_4_in_translator:uav_writedata
	wire   [27:0] fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_address;                           // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage1_to_4_in_translator:uav_address
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_write;                             // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage1_to_4_in_translator:uav_write
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_lock;                              // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage1_to_4_in_translator:uav_lock
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_read;                              // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage1_to_4_in_translator:uav_read
	wire   [31:0] fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdata;                          // fifo_stage1_to_4_in_translator:uav_readdata -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // fifo_stage1_to_4_in_translator:uav_readdatavalid -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage1_to_4_in_translator:uav_debugaccess
	wire    [3:0] fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage1_to_4_in_translator:uav_byteenable
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_data;                       // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // fifo_stage1_to_4_in_csr_translator:uav_waitrequest -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage1_to_4_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                     // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage1_to_4_in_csr_translator:uav_writedata
	wire   [27:0] fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                       // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage1_to_4_in_csr_translator:uav_address
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                         // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage1_to_4_in_csr_translator:uav_write
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                          // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage1_to_4_in_csr_translator:uav_lock
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                          // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage1_to_4_in_csr_translator:uav_read
	wire   [31:0] fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                      // fifo_stage1_to_4_in_csr_translator:uav_readdata -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // fifo_stage1_to_4_in_csr_translator:uav_readdatavalid -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage1_to_4_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage1_to_4_in_csr_translator:uav_byteenable
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                   // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // fifo_stage1_to_5_in_translator:uav_waitrequest -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage1_to_5_in_translator:uav_burstcount
	wire   [31:0] fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_writedata;                         // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage1_to_5_in_translator:uav_writedata
	wire   [27:0] fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_address;                           // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage1_to_5_in_translator:uav_address
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_write;                             // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage1_to_5_in_translator:uav_write
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_lock;                              // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage1_to_5_in_translator:uav_lock
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_read;                              // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage1_to_5_in_translator:uav_read
	wire   [31:0] fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdata;                          // fifo_stage1_to_5_in_translator:uav_readdata -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // fifo_stage1_to_5_in_translator:uav_readdatavalid -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage1_to_5_in_translator:uav_debugaccess
	wire    [3:0] fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage1_to_5_in_translator:uav_byteenable
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_data;                       // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // fifo_stage1_to_5_in_csr_translator:uav_waitrequest -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage1_to_5_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                     // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage1_to_5_in_csr_translator:uav_writedata
	wire   [27:0] fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                       // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage1_to_5_in_csr_translator:uav_address
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                         // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage1_to_5_in_csr_translator:uav_write
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                          // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage1_to_5_in_csr_translator:uav_lock
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                          // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage1_to_5_in_csr_translator:uav_read
	wire   [31:0] fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                      // fifo_stage1_to_5_in_csr_translator:uav_readdata -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // fifo_stage1_to_5_in_csr_translator:uav_readdatavalid -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage1_to_5_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage1_to_5_in_csr_translator:uav_byteenable
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                   // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // fifo_stage1_to_6_in_translator:uav_waitrequest -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage1_to_6_in_translator:uav_burstcount
	wire    [7:0] fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_writedata;                         // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage1_to_6_in_translator:uav_writedata
	wire   [27:0] fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_address;                           // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage1_to_6_in_translator:uav_address
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_write;                             // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage1_to_6_in_translator:uav_write
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_lock;                              // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage1_to_6_in_translator:uav_lock
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_read;                              // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage1_to_6_in_translator:uav_read
	wire    [7:0] fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdata;                          // fifo_stage1_to_6_in_translator:uav_readdata -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // fifo_stage1_to_6_in_translator:uav_readdatavalid -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage1_to_6_in_translator:uav_debugaccess
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage1_to_6_in_translator:uav_byteenable
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [80:0] fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_data;                       // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [80:0] fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // fifo_stage1_to_6_in_csr_translator:uav_waitrequest -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage1_to_6_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                     // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage1_to_6_in_csr_translator:uav_writedata
	wire   [27:0] fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                       // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage1_to_6_in_csr_translator:uav_address
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                         // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage1_to_6_in_csr_translator:uav_write
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                          // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage1_to_6_in_csr_translator:uav_lock
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                          // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage1_to_6_in_csr_translator:uav_read
	wire   [31:0] fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                      // fifo_stage1_to_6_in_csr_translator:uav_readdata -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // fifo_stage1_to_6_in_csr_translator:uav_readdatavalid -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage1_to_6_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage1_to_6_in_csr_translator:uav_byteenable
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                   // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // pll_pll_slave_translator:uav_waitrequest -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pll_pll_slave_translator:uav_burstcount
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                               // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pll_pll_slave_translator:uav_writedata
	wire   [27:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                                 // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> pll_pll_slave_translator:uav_address
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                                   // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> pll_pll_slave_translator:uav_write
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                    // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pll_pll_slave_translator:uav_lock
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                                    // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> pll_pll_slave_translator:uav_read
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                // pll_pll_slave_translator:uav_readdata -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // pll_pll_slave_translator:uav_readdatavalid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pll_pll_slave_translator:uav_debugaccess
	wire    [3:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pll_pll_slave_translator:uav_byteenable
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                             // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // instruction_mem_5_s1_translator:uav_waitrequest -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> instruction_mem_5_s1_translator:uav_burstcount
	wire   [31:0] instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> instruction_mem_5_s1_translator:uav_writedata
	wire   [27:0] instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_address -> instruction_mem_5_s1_translator:uav_address
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_write -> instruction_mem_5_s1_translator:uav_write
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> instruction_mem_5_s1_translator:uav_lock
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_read -> instruction_mem_5_s1_translator:uav_read
	wire   [31:0] instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // instruction_mem_5_s1_translator:uav_readdata -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // instruction_mem_5_s1_translator:uav_readdatavalid -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> instruction_mem_5_s1_translator:uav_debugaccess
	wire    [3:0] instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> instruction_mem_5_s1_translator:uav_byteenable
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_5_jtag_debug_module_translator:uav_waitrequest -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_5_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_5_jtag_debug_module_translator:uav_writedata
	wire   [27:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_5_jtag_debug_module_translator:uav_address
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_5_jtag_debug_module_translator:uav_write
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_5_jtag_debug_module_translator:uav_lock
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_5_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_5_jtag_debug_module_translator:uav_readdata -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_5_jtag_debug_module_translator:uav_readdatavalid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_5_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_5_jtag_debug_module_translator:uav_byteenable
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_5_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_5_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_5_avalon_jtag_slave_translator:uav_writedata
	wire   [27:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_5_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_5_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_5_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_5_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_5_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_5_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_5_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_5_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_5_s1_translator:uav_waitrequest -> timer_5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_5_s1_translator:uav_burstcount
	wire   [31:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_5_s1_translator:uav_writedata
	wire   [27:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_5_s1_translator:uav_address
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_5_s1_translator:uav_write
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_5_s1_translator:uav_lock
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_5_s1_translator:uav_read
	wire   [31:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_5_s1_translator:uav_readdata -> timer_5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_5_s1_translator:uav_readdatavalid -> timer_5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_5_s1_translator:uav_debugaccess
	wire    [3:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_5_s1_translator:uav_byteenable
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // fifo_stage1_to_6_out_translator:uav_waitrequest -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage1_to_6_out_translator:uav_burstcount
	wire    [7:0] fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_writedata;                        // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage1_to_6_out_translator:uav_writedata
	wire   [27:0] fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_address;                          // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage1_to_6_out_translator:uav_address
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_write;                            // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage1_to_6_out_translator:uav_write
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_lock;                             // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage1_to_6_out_translator:uav_lock
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_read;                             // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage1_to_6_out_translator:uav_read
	wire    [7:0] fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdata;                         // fifo_stage1_to_6_out_translator:uav_readdata -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // fifo_stage1_to_6_out_translator:uav_readdatavalid -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage1_to_6_out_translator:uav_debugaccess
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage1_to_6_out_translator:uav_byteenable
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [80:0] fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_data;                      // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [80:0] fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // fifo_stage5_to_6_out_translator:uav_waitrequest -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage5_to_6_out_translator:uav_burstcount
	wire   [31:0] fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_writedata;                        // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage5_to_6_out_translator:uav_writedata
	wire   [27:0] fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_address;                          // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage5_to_6_out_translator:uav_address
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_write;                            // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage5_to_6_out_translator:uav_write
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_lock;                             // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage5_to_6_out_translator:uav_lock
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_read;                             // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage5_to_6_out_translator:uav_read
	wire   [31:0] fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdata;                         // fifo_stage5_to_6_out_translator:uav_readdata -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // fifo_stage5_to_6_out_translator:uav_readdatavalid -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage5_to_6_out_translator:uav_debugaccess
	wire    [3:0] fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage5_to_6_out_translator:uav_byteenable
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_data;                      // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // fifo_stage5_to_6_in_csr_translator:uav_waitrequest -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage5_to_6_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                     // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage5_to_6_in_csr_translator:uav_writedata
	wire   [27:0] fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                       // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage5_to_6_in_csr_translator:uav_address
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                         // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage5_to_6_in_csr_translator:uav_write
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                          // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage5_to_6_in_csr_translator:uav_lock
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                          // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage5_to_6_in_csr_translator:uav_read
	wire   [31:0] fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                      // fifo_stage5_to_6_in_csr_translator:uav_readdata -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // fifo_stage5_to_6_in_csr_translator:uav_readdatavalid -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage5_to_6_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage5_to_6_in_csr_translator:uav_byteenable
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                   // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // fifo_stage4_to_5_in_csr_translator:uav_waitrequest -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage4_to_5_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                     // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage4_to_5_in_csr_translator:uav_writedata
	wire   [27:0] fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                       // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage4_to_5_in_csr_translator:uav_address
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                         // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage4_to_5_in_csr_translator:uav_write
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                          // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage4_to_5_in_csr_translator:uav_lock
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                          // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage4_to_5_in_csr_translator:uav_read
	wire   [31:0] fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                      // fifo_stage4_to_5_in_csr_translator:uav_readdata -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // fifo_stage4_to_5_in_csr_translator:uav_readdatavalid -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage4_to_5_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage4_to_5_in_csr_translator:uav_byteenable
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                   // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // instruction_mem_4_s1_translator:uav_waitrequest -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> instruction_mem_4_s1_translator:uav_burstcount
	wire   [31:0] instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> instruction_mem_4_s1_translator:uav_writedata
	wire   [27:0] instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> instruction_mem_4_s1_translator:uav_address
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> instruction_mem_4_s1_translator:uav_write
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> instruction_mem_4_s1_translator:uav_lock
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> instruction_mem_4_s1_translator:uav_read
	wire   [31:0] instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // instruction_mem_4_s1_translator:uav_readdata -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // instruction_mem_4_s1_translator:uav_readdatavalid -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> instruction_mem_4_s1_translator:uav_debugaccess
	wire    [3:0] instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> instruction_mem_4_s1_translator:uav_byteenable
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_4_jtag_debug_module_translator:uav_waitrequest -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_4_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_4_jtag_debug_module_translator:uav_writedata
	wire   [27:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_4_jtag_debug_module_translator:uav_address
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_4_jtag_debug_module_translator:uav_write
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_4_jtag_debug_module_translator:uav_lock
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_4_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_4_jtag_debug_module_translator:uav_readdata -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_4_jtag_debug_module_translator:uav_readdatavalid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_4_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_4_jtag_debug_module_translator:uav_byteenable
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_4_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_4_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_4_avalon_jtag_slave_translator:uav_writedata
	wire   [27:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_4_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_4_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_4_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_4_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_4_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_4_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_4_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_4_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_4_s1_translator:uav_waitrequest -> timer_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_4_s1_translator:uav_burstcount
	wire   [31:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_4_s1_translator:uav_writedata
	wire   [27:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_4_s1_translator:uav_address
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_4_s1_translator:uav_write
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_4_s1_translator:uav_lock
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_4_s1_translator:uav_read
	wire   [31:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_4_s1_translator:uav_readdata -> timer_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_4_s1_translator:uav_readdatavalid -> timer_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_4_s1_translator:uav_debugaccess
	wire    [3:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_4_s1_translator:uav_byteenable
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // fifo_stage1_to_5_out_translator:uav_waitrequest -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage1_to_5_out_translator:uav_burstcount
	wire   [31:0] fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_writedata;                        // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage1_to_5_out_translator:uav_writedata
	wire   [27:0] fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_address;                          // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage1_to_5_out_translator:uav_address
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_write;                            // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage1_to_5_out_translator:uav_write
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_lock;                             // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage1_to_5_out_translator:uav_lock
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_read;                             // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage1_to_5_out_translator:uav_read
	wire   [31:0] fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdata;                         // fifo_stage1_to_5_out_translator:uav_readdata -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // fifo_stage1_to_5_out_translator:uav_readdatavalid -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage1_to_5_out_translator:uav_debugaccess
	wire    [3:0] fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage1_to_5_out_translator:uav_byteenable
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_data;                      // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // fifo_stage4_to_5_out_translator:uav_waitrequest -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage4_to_5_out_translator:uav_burstcount
	wire   [31:0] fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_writedata;                        // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage4_to_5_out_translator:uav_writedata
	wire   [27:0] fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_address;                          // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage4_to_5_out_translator:uav_address
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_write;                            // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage4_to_5_out_translator:uav_write
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_lock;                             // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage4_to_5_out_translator:uav_lock
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_read;                             // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage4_to_5_out_translator:uav_read
	wire   [31:0] fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdata;                         // fifo_stage4_to_5_out_translator:uav_readdata -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // fifo_stage4_to_5_out_translator:uav_readdatavalid -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage4_to_5_out_translator:uav_debugaccess
	wire    [3:0] fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage4_to_5_out_translator:uav_byteenable
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_data;                      // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // fifo_stage5_to_6_in_translator:uav_waitrequest -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage5_to_6_in_translator:uav_burstcount
	wire   [31:0] fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_writedata;                         // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage5_to_6_in_translator:uav_writedata
	wire   [27:0] fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_address;                           // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage5_to_6_in_translator:uav_address
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_write;                             // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage5_to_6_in_translator:uav_write
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_lock;                              // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage5_to_6_in_translator:uav_lock
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_read;                              // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage5_to_6_in_translator:uav_read
	wire   [31:0] fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdata;                          // fifo_stage5_to_6_in_translator:uav_readdata -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // fifo_stage5_to_6_in_translator:uav_readdatavalid -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage5_to_6_in_translator:uav_debugaccess
	wire    [3:0] fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage5_to_6_in_translator:uav_byteenable
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_data;                       // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // instruction_mem_1_s1_translator:uav_waitrequest -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> instruction_mem_1_s1_translator:uav_burstcount
	wire   [31:0] instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> instruction_mem_1_s1_translator:uav_writedata
	wire   [27:0] instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> instruction_mem_1_s1_translator:uav_address
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> instruction_mem_1_s1_translator:uav_write
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> instruction_mem_1_s1_translator:uav_lock
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> instruction_mem_1_s1_translator:uav_read
	wire   [31:0] instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // instruction_mem_1_s1_translator:uav_readdata -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // instruction_mem_1_s1_translator:uav_readdatavalid -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> instruction_mem_1_s1_translator:uav_debugaccess
	wire    [3:0] instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> instruction_mem_1_s1_translator:uav_byteenable
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_1_jtag_debug_module_translator:uav_waitrequest -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_1_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_1_jtag_debug_module_translator:uav_writedata
	wire   [27:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_1_jtag_debug_module_translator:uav_address
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_1_jtag_debug_module_translator:uav_write
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_1_jtag_debug_module_translator:uav_lock
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_1_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_1_jtag_debug_module_translator:uav_readdata -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_1_jtag_debug_module_translator:uav_readdatavalid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_1_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_1_jtag_debug_module_translator:uav_byteenable
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_1_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_1_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_1_avalon_jtag_slave_translator:uav_writedata
	wire   [27:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_1_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_1_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_1_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_1_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_1_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_1_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_1_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_1_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	wire   [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	wire   [27:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	wire   [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	wire    [3:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // fifo_0_stage1_to_2_out_translator:uav_waitrequest -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_stage1_to_2_out_translator:uav_burstcount
	wire   [31:0] fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata;                      // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_stage1_to_2_out_translator:uav_writedata
	wire   [27:0] fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address;                        // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_stage1_to_2_out_translator:uav_address
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write;                          // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_stage1_to_2_out_translator:uav_write
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock;                           // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_stage1_to_2_out_translator:uav_lock
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read;                           // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_stage1_to_2_out_translator:uav_read
	wire   [31:0] fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata;                       // fifo_0_stage1_to_2_out_translator:uav_readdata -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // fifo_0_stage1_to_2_out_translator:uav_readdatavalid -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_stage1_to_2_out_translator:uav_debugaccess
	wire    [3:0] fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_stage1_to_2_out_translator:uav_byteenable
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data;                    // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // fifo_1_stage1_to_2_out_translator:uav_waitrequest -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_stage1_to_2_out_translator:uav_burstcount
	wire   [31:0] fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata;                      // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_stage1_to_2_out_translator:uav_writedata
	wire   [27:0] fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address;                        // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_stage1_to_2_out_translator:uav_address
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write;                          // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_stage1_to_2_out_translator:uav_write
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock;                           // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_stage1_to_2_out_translator:uav_lock
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read;                           // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_stage1_to_2_out_translator:uav_read
	wire   [31:0] fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata;                       // fifo_1_stage1_to_2_out_translator:uav_readdata -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // fifo_1_stage1_to_2_out_translator:uav_readdatavalid -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_stage1_to_2_out_translator:uav_debugaccess
	wire    [3:0] fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_stage1_to_2_out_translator:uav_byteenable
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data;                    // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // fifo_2_stage1_to_2_out_translator:uav_waitrequest -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_stage1_to_2_out_translator:uav_burstcount
	wire   [31:0] fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata;                      // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_stage1_to_2_out_translator:uav_writedata
	wire   [27:0] fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address;                        // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_stage1_to_2_out_translator:uav_address
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write;                          // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_stage1_to_2_out_translator:uav_write
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock;                           // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_stage1_to_2_out_translator:uav_lock
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read;                           // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_stage1_to_2_out_translator:uav_read
	wire   [31:0] fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata;                       // fifo_2_stage1_to_2_out_translator:uav_readdata -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // fifo_2_stage1_to_2_out_translator:uav_readdatavalid -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_stage1_to_2_out_translator:uav_debugaccess
	wire    [3:0] fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_stage1_to_2_out_translator:uav_byteenable
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data;                    // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // fifo_stage2_to_3_in_translator:uav_waitrequest -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage2_to_3_in_translator:uav_burstcount
	wire   [31:0] fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_writedata;                         // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage2_to_3_in_translator:uav_writedata
	wire   [27:0] fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_address;                           // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage2_to_3_in_translator:uav_address
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_write;                             // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage2_to_3_in_translator:uav_write
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_lock;                              // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage2_to_3_in_translator:uav_lock
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_read;                              // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage2_to_3_in_translator:uav_read
	wire   [31:0] fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_readdata;                          // fifo_stage2_to_3_in_translator:uav_readdata -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // fifo_stage2_to_3_in_translator:uav_readdatavalid -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage2_to_3_in_translator:uav_debugaccess
	wire    [3:0] fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage2_to_3_in_translator:uav_byteenable
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_data;                       // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // fifo_stage2_to_3_in_csr_translator:uav_waitrequest -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage2_to_3_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                     // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage2_to_3_in_csr_translator:uav_writedata
	wire   [27:0] fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                       // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage2_to_3_in_csr_translator:uav_address
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                         // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage2_to_3_in_csr_translator:uav_write
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                          // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage2_to_3_in_csr_translator:uav_lock
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                          // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage2_to_3_in_csr_translator:uav_read
	wire   [31:0] fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                      // fifo_stage2_to_3_in_csr_translator:uav_readdata -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // fifo_stage2_to_3_in_csr_translator:uav_readdatavalid -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage2_to_3_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage2_to_3_in_csr_translator:uav_byteenable
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                   // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // instruction_mem_2_s1_translator:uav_waitrequest -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> instruction_mem_2_s1_translator:uav_burstcount
	wire   [31:0] instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> instruction_mem_2_s1_translator:uav_writedata
	wire   [27:0] instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> instruction_mem_2_s1_translator:uav_address
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> instruction_mem_2_s1_translator:uav_write
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> instruction_mem_2_s1_translator:uav_lock
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> instruction_mem_2_s1_translator:uav_read
	wire   [31:0] instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // instruction_mem_2_s1_translator:uav_readdata -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // instruction_mem_2_s1_translator:uav_readdatavalid -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> instruction_mem_2_s1_translator:uav_debugaccess
	wire    [3:0] instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> instruction_mem_2_s1_translator:uav_byteenable
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_2_jtag_debug_module_translator:uav_waitrequest -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_2_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_2_jtag_debug_module_translator:uav_writedata
	wire   [27:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_2_jtag_debug_module_translator:uav_address
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_2_jtag_debug_module_translator:uav_write
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_2_jtag_debug_module_translator:uav_lock
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_2_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_2_jtag_debug_module_translator:uav_readdata -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_2_jtag_debug_module_translator:uav_readdatavalid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_2_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_2_jtag_debug_module_translator:uav_byteenable
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_2_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_2_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_2_avalon_jtag_slave_translator:uav_writedata
	wire   [27:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_2_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_2_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_2_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_2_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_2_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_2_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_2_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_2_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_2_s1_translator:uav_waitrequest -> timer_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_2_s1_translator:uav_burstcount
	wire   [31:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_2_s1_translator:uav_writedata
	wire   [27:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_2_s1_translator:uav_address
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_2_s1_translator:uav_write
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_2_s1_translator:uav_lock
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_2_s1_translator:uav_read
	wire   [31:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_2_s1_translator:uav_readdata -> timer_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_2_s1_translator:uav_readdatavalid -> timer_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_2_s1_translator:uav_debugaccess
	wire    [3:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_2_s1_translator:uav_byteenable
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // fifo_stage2_to_3_out_translator:uav_waitrequest -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage2_to_3_out_translator:uav_burstcount
	wire   [31:0] fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_writedata;                        // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage2_to_3_out_translator:uav_writedata
	wire   [27:0] fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_address;                          // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage2_to_3_out_translator:uav_address
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_write;                            // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage2_to_3_out_translator:uav_write
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_lock;                             // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage2_to_3_out_translator:uav_lock
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_read;                             // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage2_to_3_out_translator:uav_read
	wire   [31:0] fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_readdata;                         // fifo_stage2_to_3_out_translator:uav_readdata -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // fifo_stage2_to_3_out_translator:uav_readdatavalid -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage2_to_3_out_translator:uav_debugaccess
	wire    [3:0] fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage2_to_3_out_translator:uav_byteenable
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_data;                      // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // fifo_stage3_to_4_in_translator:uav_waitrequest -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage3_to_4_in_translator:uav_burstcount
	wire   [31:0] fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_writedata;                         // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage3_to_4_in_translator:uav_writedata
	wire   [27:0] fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_address;                           // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage3_to_4_in_translator:uav_address
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_write;                             // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage3_to_4_in_translator:uav_write
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_lock;                              // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage3_to_4_in_translator:uav_lock
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_read;                              // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage3_to_4_in_translator:uav_read
	wire   [31:0] fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdata;                          // fifo_stage3_to_4_in_translator:uav_readdata -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // fifo_stage3_to_4_in_translator:uav_readdatavalid -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage3_to_4_in_translator:uav_debugaccess
	wire    [3:0] fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage3_to_4_in_translator:uav_byteenable
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_data;                       // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // fifo_stage3_to_4_in_csr_translator:uav_waitrequest -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage3_to_4_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                     // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage3_to_4_in_csr_translator:uav_writedata
	wire   [27:0] fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                       // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage3_to_4_in_csr_translator:uav_address
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                         // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage3_to_4_in_csr_translator:uav_write
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                          // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage3_to_4_in_csr_translator:uav_lock
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                          // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage3_to_4_in_csr_translator:uav_read
	wire   [31:0] fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                      // fifo_stage3_to_4_in_csr_translator:uav_readdata -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // fifo_stage3_to_4_in_csr_translator:uav_readdatavalid -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage3_to_4_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage3_to_4_in_csr_translator:uav_byteenable
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                   // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // instruction_mem_3_s1_translator:uav_waitrequest -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> instruction_mem_3_s1_translator:uav_burstcount
	wire   [31:0] instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> instruction_mem_3_s1_translator:uav_writedata
	wire   [27:0] instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> instruction_mem_3_s1_translator:uav_address
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> instruction_mem_3_s1_translator:uav_write
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> instruction_mem_3_s1_translator:uav_lock
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> instruction_mem_3_s1_translator:uav_read
	wire   [31:0] instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // instruction_mem_3_s1_translator:uav_readdata -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // instruction_mem_3_s1_translator:uav_readdatavalid -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> instruction_mem_3_s1_translator:uav_debugaccess
	wire    [3:0] instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> instruction_mem_3_s1_translator:uav_byteenable
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_3_jtag_debug_module_translator:uav_waitrequest -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_3_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_3_jtag_debug_module_translator:uav_writedata
	wire   [27:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_3_jtag_debug_module_translator:uav_address
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_3_jtag_debug_module_translator:uav_write
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_3_jtag_debug_module_translator:uav_lock
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_3_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_3_jtag_debug_module_translator:uav_readdata -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_3_jtag_debug_module_translator:uav_readdatavalid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_3_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_3_jtag_debug_module_translator:uav_byteenable
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_3_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_3_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_3_avalon_jtag_slave_translator:uav_writedata
	wire   [27:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_3_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_3_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_3_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_3_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_3_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_3_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_3_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_3_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_3_s1_translator:uav_waitrequest -> timer_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_3_s1_translator:uav_burstcount
	wire   [31:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_3_s1_translator:uav_writedata
	wire   [27:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_3_s1_translator:uav_address
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_3_s1_translator:uav_write
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_3_s1_translator:uav_lock
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_3_s1_translator:uav_read
	wire   [31:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_3_s1_translator:uav_readdata -> timer_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_3_s1_translator:uav_readdatavalid -> timer_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_3_s1_translator:uav_debugaccess
	wire    [3:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_3_s1_translator:uav_byteenable
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // fifo_stage1_to_4_out_translator:uav_waitrequest -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage1_to_4_out_translator:uav_burstcount
	wire   [31:0] fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_writedata;                        // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage1_to_4_out_translator:uav_writedata
	wire   [27:0] fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_address;                          // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage1_to_4_out_translator:uav_address
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_write;                            // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage1_to_4_out_translator:uav_write
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_lock;                             // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage1_to_4_out_translator:uav_lock
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_read;                             // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage1_to_4_out_translator:uav_read
	wire   [31:0] fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdata;                         // fifo_stage1_to_4_out_translator:uav_readdata -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // fifo_stage1_to_4_out_translator:uav_readdatavalid -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage1_to_4_out_translator:uav_debugaccess
	wire    [3:0] fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage1_to_4_out_translator:uav_byteenable
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_data;                      // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // fifo_stage3_to_4_out_translator:uav_waitrequest -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage3_to_4_out_translator:uav_burstcount
	wire   [31:0] fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_writedata;                        // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage3_to_4_out_translator:uav_writedata
	wire   [27:0] fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_address;                          // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage3_to_4_out_translator:uav_address
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_write;                            // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage3_to_4_out_translator:uav_write
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_lock;                             // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage3_to_4_out_translator:uav_lock
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_read;                             // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage3_to_4_out_translator:uav_read
	wire   [31:0] fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdata;                         // fifo_stage3_to_4_out_translator:uav_readdata -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // fifo_stage3_to_4_out_translator:uav_readdatavalid -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage3_to_4_out_translator:uav_debugaccess
	wire    [3:0] fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage3_to_4_out_translator:uav_byteenable
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_data;                      // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // fifo_stage4_to_5_in_translator:uav_waitrequest -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_stage4_to_5_in_translator:uav_burstcount
	wire   [31:0] fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_writedata;                         // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_stage4_to_5_in_translator:uav_writedata
	wire   [27:0] fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_address;                           // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_stage4_to_5_in_translator:uav_address
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_write;                             // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_stage4_to_5_in_translator:uav_write
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_lock;                              // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_stage4_to_5_in_translator:uav_lock
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_read;                              // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_stage4_to_5_in_translator:uav_read
	wire   [31:0] fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdata;                          // fifo_stage4_to_5_in_translator:uav_readdata -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // fifo_stage4_to_5_in_translator:uav_readdatavalid -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_stage4_to_5_in_translator:uav_debugaccess
	wire    [3:0] fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_stage4_to_5_in_translator:uav_byteenable
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_data;                       // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [106:0] cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router:sink_ready -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [106:0] cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_001:sink_ready -> cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [106:0] cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_002:sink_ready -> cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [106:0] cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_003:sink_ready -> cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [106:0] cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_004:sink_ready -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [106:0] cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_005:sink_ready -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire          cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire          cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire  [106:0] cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire          cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_006:sink_ready -> cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	wire          cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	wire          cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	wire  [106:0] cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	wire          cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_007:sink_ready -> cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_008:sink_endofpacket
	wire          cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_008:sink_valid
	wire          cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_008:sink_startofpacket
	wire  [106:0] cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_008:sink_data
	wire          cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_008:sink_ready -> cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_009:sink_endofpacket
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_009:sink_valid
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_009:sink_startofpacket
	wire  [106:0] cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_009:sink_data
	wire          cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_009:sink_ready -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_010:sink_endofpacket
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_010:sink_valid
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_010:sink_startofpacket
	wire  [106:0] cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_010:sink_data
	wire          cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_010:sink_ready -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_011:sink_endofpacket
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_011:sink_valid
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_011:sink_startofpacket
	wire  [106:0] cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_011:sink_data
	wire          cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_011:sink_ready -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [106:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router:sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [106:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_001:sink_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [106:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_002:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [106:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid;                           // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [106:0] fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data;                            // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_004:sink_ready -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                       // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [106:0] fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                        // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_005:sink_ready -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid;                           // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [106:0] fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data;                            // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_006:sink_ready -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid;                           // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [106:0] fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data;                            // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_007:sink_ready -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                       // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [106:0] fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                        // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_008:sink_ready -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                       // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [106:0] fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                        // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_009:sink_ready -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_valid;                             // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [106:0] fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_data;                              // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_010:sink_ready -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                         // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [106:0] fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                          // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_011:sink_ready -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_valid;                             // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [106:0] fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_data;                              // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_012:sink_ready -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                         // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [106:0] fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                          // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_013:sink_ready -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_valid;                             // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire   [79:0] fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_data;                              // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_014:sink_ready -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                         // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [106:0] fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                          // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_015:sink_ready -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                   // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [106:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                                    // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_016:sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [106:0] instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_017:sink_ready -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [106:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_018:sink_ready -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [106:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_019:sink_ready -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [106:0] timer_5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          timer_5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_020:sink_ready -> timer_5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_valid;                            // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire   [79:0] fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_data;                             // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire          fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_021:sink_ready -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_valid;                            // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [106:0] fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_data;                             // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire          fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_022:sink_ready -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                         // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire  [106:0] fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                          // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire          fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_023:sink_ready -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                         // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire  [106:0] fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                          // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire          fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_024:sink_ready -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire  [106:0] instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire          instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_025:sink_ready -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire  [106:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire          cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_026:sink_ready -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire  [106:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire          jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_027:sink_ready -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire  [106:0] timer_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire          timer_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_028:sink_ready -> timer_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_valid;                            // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire  [106:0] fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_data;                             // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire          fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_029:sink_ready -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_valid;                            // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire  [106:0] fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_data;                             // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire          fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_030:sink_ready -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_valid;                             // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	wire  [106:0] fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_data;                              // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	wire          fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_031:sink_ready -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	wire  [106:0] instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	wire          instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_032:sink_ready -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_033:sink_endofpacket
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_033:sink_valid
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_033:sink_startofpacket
	wire  [106:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_033:sink_data
	wire          cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_033:sink_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_034:sink_endofpacket
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_034:sink_valid
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_034:sink_startofpacket
	wire  [106:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_034:sink_data
	wire          jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_034:sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_035:sink_endofpacket
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_035:sink_valid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_035:sink_startofpacket
	wire  [106:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_035:sink_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_035:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_036:sink_endofpacket
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid;                          // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_036:sink_valid
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_036:sink_startofpacket
	wire  [106:0] fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data;                           // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_036:sink_data
	wire          fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_036:sink_ready -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_037:sink_endofpacket
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid;                          // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_037:sink_valid
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_037:sink_startofpacket
	wire  [106:0] fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data;                           // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_037:sink_data
	wire          fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_037:sink_ready -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_038:sink_endofpacket
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid;                          // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_038:sink_valid
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_038:sink_startofpacket
	wire  [106:0] fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data;                           // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_038:sink_data
	wire          fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_038:sink_ready -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_039:sink_endofpacket
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_valid;                             // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_039:sink_valid
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_039:sink_startofpacket
	wire  [106:0] fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_data;                              // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_039:sink_data
	wire          fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_039:sink_ready -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_040:sink_endofpacket
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                         // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_040:sink_valid
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_040:sink_startofpacket
	wire  [106:0] fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                          // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_040:sink_data
	wire          fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_040:sink_ready -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_041:sink_endofpacket
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_041:sink_valid
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_041:sink_startofpacket
	wire  [106:0] instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_041:sink_data
	wire          instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_041:sink_ready -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_042:sink_endofpacket
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_042:sink_valid
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_042:sink_startofpacket
	wire  [106:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_042:sink_data
	wire          cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_042:sink_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_043:sink_endofpacket
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_043:sink_valid
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_043:sink_startofpacket
	wire  [106:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_043:sink_data
	wire          jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_043:sink_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_044:sink_endofpacket
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_044:sink_valid
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_044:sink_startofpacket
	wire  [106:0] timer_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_044:sink_data
	wire          timer_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_044:sink_ready -> timer_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_045:sink_endofpacket
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_valid;                            // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_045:sink_valid
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_045:sink_startofpacket
	wire  [106:0] fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_data;                             // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_045:sink_data
	wire          fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_045:sink_ready -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_046:sink_endofpacket
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_valid;                             // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_046:sink_valid
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_046:sink_startofpacket
	wire  [106:0] fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_data;                              // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_046:sink_data
	wire          fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_046:sink_ready -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_047:sink_endofpacket
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                         // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_047:sink_valid
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_047:sink_startofpacket
	wire  [106:0] fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                          // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_047:sink_data
	wire          fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_047:sink_ready -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_048:sink_endofpacket
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_048:sink_valid
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_048:sink_startofpacket
	wire  [106:0] instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_048:sink_data
	wire          instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_048:sink_ready -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_049:sink_endofpacket
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_049:sink_valid
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_049:sink_startofpacket
	wire  [106:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_049:sink_data
	wire          cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_049:sink_ready -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_050:sink_endofpacket
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_050:sink_valid
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_050:sink_startofpacket
	wire  [106:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_050:sink_data
	wire          jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_050:sink_ready -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_051:sink_endofpacket
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_051:sink_valid
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_051:sink_startofpacket
	wire  [106:0] timer_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_051:sink_data
	wire          timer_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_051:sink_ready -> timer_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_052:sink_endofpacket
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_valid;                            // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_052:sink_valid
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_052:sink_startofpacket
	wire  [106:0] fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_data;                             // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_052:sink_data
	wire          fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_052:sink_ready -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_053:sink_endofpacket
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_valid;                            // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_053:sink_valid
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_053:sink_startofpacket
	wire  [106:0] fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_data;                             // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_053:sink_data
	wire          fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_053:sink_ready -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_054:sink_endofpacket
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_valid;                             // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_054:sink_valid
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_054:sink_startofpacket
	wire  [106:0] fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_data;                              // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_054:sink_data
	wire          fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_054:sink_ready -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                        // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                              // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                      // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [106:0] addr_router_src_data;                                                                               // addr_router:src_data -> limiter:cmd_sink_data
	wire   [54:0] addr_router_src_channel;                                                                            // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                              // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                        // limiter:rsp_src_endofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                              // limiter:rsp_src_valid -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                      // limiter:rsp_src_startofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_rsp_src_data;                                                                               // limiter:rsp_src_data -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] limiter_rsp_src_channel;                                                                            // limiter:rsp_src_channel -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                              // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_004_src_endofpacket;                                                                    // addr_router_004:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_004_src_valid;                                                                          // addr_router_004:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_004_src_startofpacket;                                                                  // addr_router_004:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [106:0] addr_router_004_src_data;                                                                           // addr_router_004:src_data -> limiter_001:cmd_sink_data
	wire   [54:0] addr_router_004_src_channel;                                                                        // addr_router_004:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_004_src_ready;                                                                          // limiter_001:cmd_sink_ready -> addr_router_004:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                    // limiter_001:rsp_src_endofpacket -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                          // limiter_001:rsp_src_valid -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                  // limiter_001:rsp_src_startofpacket -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_001_rsp_src_data;                                                                           // limiter_001:rsp_src_data -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] limiter_001_rsp_src_channel;                                                                        // limiter_001:rsp_src_channel -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                          // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_005_src_endofpacket;                                                                    // addr_router_005:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_005_src_valid;                                                                          // addr_router_005:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_005_src_startofpacket;                                                                  // addr_router_005:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire  [106:0] addr_router_005_src_data;                                                                           // addr_router_005:src_data -> limiter_002:cmd_sink_data
	wire   [54:0] addr_router_005_src_channel;                                                                        // addr_router_005:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_005_src_ready;                                                                          // limiter_002:cmd_sink_ready -> addr_router_005:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                    // limiter_002:rsp_src_endofpacket -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                          // limiter_002:rsp_src_valid -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                  // limiter_002:rsp_src_startofpacket -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_002_rsp_src_data;                                                                           // limiter_002:rsp_src_data -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] limiter_002_rsp_src_channel;                                                                        // limiter_002:rsp_src_channel -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_002_rsp_src_ready;                                                                          // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire          addr_router_009_src_endofpacket;                                                                    // addr_router_009:src_endofpacket -> limiter_003:cmd_sink_endofpacket
	wire          addr_router_009_src_valid;                                                                          // addr_router_009:src_valid -> limiter_003:cmd_sink_valid
	wire          addr_router_009_src_startofpacket;                                                                  // addr_router_009:src_startofpacket -> limiter_003:cmd_sink_startofpacket
	wire  [106:0] addr_router_009_src_data;                                                                           // addr_router_009:src_data -> limiter_003:cmd_sink_data
	wire   [54:0] addr_router_009_src_channel;                                                                        // addr_router_009:src_channel -> limiter_003:cmd_sink_channel
	wire          addr_router_009_src_ready;                                                                          // limiter_003:cmd_sink_ready -> addr_router_009:src_ready
	wire          limiter_003_rsp_src_endofpacket;                                                                    // limiter_003:rsp_src_endofpacket -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_003_rsp_src_valid;                                                                          // limiter_003:rsp_src_valid -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_003_rsp_src_startofpacket;                                                                  // limiter_003:rsp_src_startofpacket -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_003_rsp_src_data;                                                                           // limiter_003:rsp_src_data -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] limiter_003_rsp_src_channel;                                                                        // limiter_003:rsp_src_channel -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_003_rsp_src_ready;                                                                          // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_003:rsp_src_ready
	wire          addr_router_010_src_endofpacket;                                                                    // addr_router_010:src_endofpacket -> limiter_004:cmd_sink_endofpacket
	wire          addr_router_010_src_valid;                                                                          // addr_router_010:src_valid -> limiter_004:cmd_sink_valid
	wire          addr_router_010_src_startofpacket;                                                                  // addr_router_010:src_startofpacket -> limiter_004:cmd_sink_startofpacket
	wire  [106:0] addr_router_010_src_data;                                                                           // addr_router_010:src_data -> limiter_004:cmd_sink_data
	wire   [54:0] addr_router_010_src_channel;                                                                        // addr_router_010:src_channel -> limiter_004:cmd_sink_channel
	wire          addr_router_010_src_ready;                                                                          // limiter_004:cmd_sink_ready -> addr_router_010:src_ready
	wire          limiter_004_rsp_src_endofpacket;                                                                    // limiter_004:rsp_src_endofpacket -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_004_rsp_src_valid;                                                                          // limiter_004:rsp_src_valid -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_004_rsp_src_startofpacket;                                                                  // limiter_004:rsp_src_startofpacket -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_004_rsp_src_data;                                                                           // limiter_004:rsp_src_data -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] limiter_004_rsp_src_channel;                                                                        // limiter_004:rsp_src_channel -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_004_rsp_src_ready;                                                                          // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_004:rsp_src_ready
	wire          addr_router_011_src_endofpacket;                                                                    // addr_router_011:src_endofpacket -> limiter_005:cmd_sink_endofpacket
	wire          addr_router_011_src_valid;                                                                          // addr_router_011:src_valid -> limiter_005:cmd_sink_valid
	wire          addr_router_011_src_startofpacket;                                                                  // addr_router_011:src_startofpacket -> limiter_005:cmd_sink_startofpacket
	wire  [106:0] addr_router_011_src_data;                                                                           // addr_router_011:src_data -> limiter_005:cmd_sink_data
	wire   [54:0] addr_router_011_src_channel;                                                                        // addr_router_011:src_channel -> limiter_005:cmd_sink_channel
	wire          addr_router_011_src_ready;                                                                          // limiter_005:cmd_sink_ready -> addr_router_011:src_ready
	wire          limiter_005_rsp_src_endofpacket;                                                                    // limiter_005:rsp_src_endofpacket -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_005_rsp_src_valid;                                                                          // limiter_005:rsp_src_valid -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_005_rsp_src_startofpacket;                                                                  // limiter_005:rsp_src_startofpacket -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_005_rsp_src_data;                                                                           // limiter_005:rsp_src_data -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] limiter_005_rsp_src_channel;                                                                        // limiter_005:rsp_src_channel -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_005_rsp_src_ready;                                                                          // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_005:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                  // burst_adapter:source0_endofpacket -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                        // burst_adapter:source0_valid -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                // burst_adapter:source0_startofpacket -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [79:0] burst_adapter_source0_data;                                                                         // burst_adapter:source0_data -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                        // fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [54:0] burst_adapter_source0_channel;                                                                      // burst_adapter:source0_channel -> fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                              // burst_adapter_001:source0_endofpacket -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                    // burst_adapter_001:source0_valid -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                            // burst_adapter_001:source0_startofpacket -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [79:0] burst_adapter_001_source0_data;                                                                     // burst_adapter_001:source0_data -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                    // fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [54:0] burst_adapter_001_source0_channel;                                                                  // burst_adapter_001:source0_channel -> fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                     // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, addr_router_005:reset, addr_router_006:reset, addr_router_007:reset, addr_router_008:reset, addr_router_009:reset, addr_router_010:reset, addr_router_011:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_demux_006:reset, cmd_xbar_demux_007:reset, cmd_xbar_demux_008:reset, cmd_xbar_demux_009:reset, cmd_xbar_demux_010:reset, cmd_xbar_demux_011:reset, cmd_xbar_mux:reset, cmd_xbar_mux_018:reset, cmd_xbar_mux_026:reset, cmd_xbar_mux_033:reset, cmd_xbar_mux_042:reset, cmd_xbar_mux_049:reset, cpu_0:reset_n, cpu_0_data_master_translator:reset, cpu_0_data_master_translator_avalon_universal_master_0_agent:reset, cpu_0_instruction_master_translator:reset, cpu_0_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_0_jtag_debug_module_translator:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_1:reset_n, cpu_1_data_master_translator:reset, cpu_1_data_master_translator_avalon_universal_master_0_agent:reset, cpu_1_instruction_master_translator:reset, cpu_1_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_1_jtag_debug_module_translator:reset, cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_2:reset_n, cpu_2_data_master_translator:reset, cpu_2_data_master_translator_avalon_universal_master_0_agent:reset, cpu_2_instruction_master_translator:reset, cpu_2_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_2_jtag_debug_module_translator:reset, cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_3:reset_n, cpu_3_data_master_translator:reset, cpu_3_data_master_translator_avalon_universal_master_0_agent:reset, cpu_3_instruction_master_translator:reset, cpu_3_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_3_jtag_debug_module_translator:reset, cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_4:reset_n, cpu_4_data_master_translator:reset, cpu_4_data_master_translator_avalon_universal_master_0_agent:reset, cpu_4_instruction_master_translator:reset, cpu_4_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_4_jtag_debug_module_translator:reset, cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_5:reset_n, cpu_5_data_master_translator:reset, cpu_5_data_master_translator_avalon_universal_master_0_agent:reset, cpu_5_instruction_master_translator:reset, cpu_5_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_5_jtag_debug_module_translator:reset, cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_018:reset, id_router_026:reset, id_router_033:reset, id_router_042:reset, id_router_049:reset, irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, irq_mapper_004:reset, irq_mapper_005:reset, limiter:reset, limiter_001:reset, limiter_002:reset, limiter_003:reset, limiter_004:reset, limiter_005:reset, rsp_xbar_demux:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_033:reset, rsp_xbar_demux_042:reset, rsp_xbar_demux_049:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, rsp_xbar_mux_003:reset, rsp_xbar_mux_004:reset, rsp_xbar_mux_005:reset, rsp_xbar_mux_006:reset, rsp_xbar_mux_007:reset, rsp_xbar_mux_008:reset, rsp_xbar_mux_009:reset, rsp_xbar_mux_010:reset, rsp_xbar_mux_011:reset]
	wire          rst_controller_001_reset_out_reset;                                                                 // rst_controller_001:reset_out -> [id_router_002:reset, id_router_003:reset, id_router_016:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pll:reset, pll_pll_slave_translator:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_016:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cpu_0_jtag_debug_module_reset_reset;                                                                // cpu_0:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in1, rst_controller_007:reset_in1, rst_controller_008:reset_in1, rst_controller_009:reset_in1, rst_controller_010:reset_in1, rst_controller_015:reset_in1]
	wire          rst_controller_002_reset_out_reset;                                                                 // rst_controller_002:reset_out -> [cmd_xbar_mux_032:reset, id_router_032:reset, id_router_034:reset, id_router_035:reset, instruction_mem_1:reset, instruction_mem_1_s1_translator:reset, instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:reset, instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, jtag_uart_1:rst_n, jtag_uart_1_avalon_jtag_slave_translator:reset, jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_032:reset, rsp_xbar_demux_034:reset, rsp_xbar_demux_035:reset, timer_1:reset_n, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cpu_1_jtag_debug_module_reset_reset;                                                                // cpu_1:jtag_debug_module_resetrequest -> [rst_controller_002:reset_in1, rst_controller_007:reset_in2, rst_controller_011:reset_in1, rst_controller_015:reset_in2]
	wire          rst_controller_003_reset_out_reset;                                                                 // rst_controller_003:reset_out -> [cmd_xbar_mux_041:reset, id_router_041:reset, id_router_044:reset, instruction_mem_2:reset, instruction_mem_2_s1_translator:reset, instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:reset, instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_041:reset, rsp_xbar_demux_044:reset, timer_2:reset_n, timer_2_s1_translator:reset, timer_2_s1_translator_avalon_universal_slave_0_agent:reset, timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_004_reset_out_reset;                                                                 // rst_controller_004:reset_out -> [cmd_xbar_mux_048:reset, id_router_048:reset, id_router_050:reset, id_router_051:reset, instruction_mem_3:reset, instruction_mem_3_s1_translator:reset, instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:reset, instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, jtag_uart_3:rst_n, jtag_uart_3_avalon_jtag_slave_translator:reset, jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_048:reset, rsp_xbar_demux_050:reset, rsp_xbar_demux_051:reset, timer_3:reset_n, timer_3_s1_translator:reset, timer_3_s1_translator_avalon_universal_slave_0_agent:reset, timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cpu_3_jtag_debug_module_reset_reset;                                                                // cpu_3:jtag_debug_module_resetrequest -> [rst_controller_004:reset_in1, rst_controller_008:reset_in2, rst_controller_012:reset_in2, rst_controller_013:reset_in1, rst_controller_015:reset_in4]
	wire          rst_controller_005_reset_out_reset;                                                                 // rst_controller_005:reset_out -> [cmd_xbar_mux_025:reset, id_router_025:reset, id_router_027:reset, id_router_028:reset, instruction_mem_4:reset, instruction_mem_4_s1_translator:reset, instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:reset, instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, jtag_uart_4:rst_n, jtag_uart_4_avalon_jtag_slave_translator:reset, jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, timer_4:reset_n, timer_4_s1_translator:reset, timer_4_s1_translator_avalon_universal_slave_0_agent:reset, timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cpu_4_jtag_debug_module_reset_reset;                                                                // cpu_4:jtag_debug_module_resetrequest -> [rst_controller_005:reset_in1, rst_controller_009:reset_in2, rst_controller_013:reset_in2, rst_controller_014:reset_in1, rst_controller_015:reset_in5]
	wire          rst_controller_006_reset_out_reset;                                                                 // rst_controller_006:reset_out -> [cmd_xbar_mux_017:reset, id_router_017:reset, id_router_019:reset, id_router_020:reset, instruction_mem_5:reset, instruction_mem_5_s1_translator:reset, instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:reset, instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, jtag_uart_5:rst_n, jtag_uart_5_avalon_jtag_slave_translator:reset, jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, timer_5:reset_n, timer_5_s1_translator:reset, timer_5_s1_translator_avalon_universal_slave_0_agent:reset, timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cpu_5_jtag_debug_module_reset_reset;                                                                // cpu_5:jtag_debug_module_resetrequest -> [rst_controller_006:reset_in1, rst_controller_010:reset_in2, rst_controller_014:reset_in2, rst_controller_015:reset_in6]
	wire          rst_controller_007_reset_out_reset;                                                                 // rst_controller_007:reset_out -> [cmd_xbar_mux_005:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, fifo_0_stage1_to_2:reset_n, fifo_0_stage1_to_2_in_csr_translator:reset, fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_stage1_to_2_in_translator:reset, fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:reset, fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_stage1_to_2_out_translator:reset, fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:reset, fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_stage1_to_2:reset_n, fifo_1_stage1_to_2_in_csr_translator:reset, fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_stage1_to_2_in_translator:reset, fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:reset, fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_stage1_to_2_out_translator:reset, fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:reset, fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_stage1_to_2:reset_n, fifo_2_stage1_to_2_in_csr_translator:reset, fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_stage1_to_2_in_translator:reset, fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:reset, fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_stage1_to_2_out_translator:reset, fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:reset, fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_036:reset, id_router_037:reset, id_router_038:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_036:reset, rsp_xbar_demux_037:reset, rsp_xbar_demux_038:reset]
	wire          rst_controller_008_reset_out_reset;                                                                 // rst_controller_008:reset_out -> [cmd_xbar_mux_011:reset, fifo_stage1_to_4:reset_n, fifo_stage1_to_4_in_csr_translator:reset, fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage1_to_4_in_translator:reset, fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:reset, fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage1_to_4_out_translator:reset, fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:reset, fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_010:reset, id_router_011:reset, id_router_052:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_052:reset]
	wire          rst_controller_009_reset_out_reset;                                                                 // rst_controller_009:reset_out -> [cmd_xbar_mux_013:reset, fifo_stage1_to_5:reset_n, fifo_stage1_to_5_in_csr_translator:reset, fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage1_to_5_in_translator:reset, fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:reset, fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage1_to_5_out_translator:reset, fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:reset, fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_012:reset, id_router_013:reset, id_router_029:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_029:reset]
	wire          rst_controller_010_reset_out_reset;                                                                 // rst_controller_010:reset_out -> [burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_mux_015:reset, fifo_stage1_to_6:reset_n, fifo_stage1_to_6_in_csr_translator:reset, fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage1_to_6_in_translator:reset, fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent:reset, fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage1_to_6_out_translator:reset, fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent:reset, fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_014:reset, id_router_015:reset, id_router_021:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_021:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_011_reset_out_reset;                                                                 // rst_controller_011:reset_out -> [cmd_xbar_mux_040:reset, fifo_stage2_to_3:reset_n, fifo_stage2_to_3_in_csr_translator:reset, fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage2_to_3_in_translator:reset, fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:reset, fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage2_to_3_out_translator:reset, fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:reset, fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_039:reset, id_router_040:reset, id_router_045:reset, rsp_xbar_demux_039:reset, rsp_xbar_demux_040:reset, rsp_xbar_demux_045:reset]
	wire          rst_controller_012_reset_out_reset;                                                                 // rst_controller_012:reset_out -> [cmd_xbar_mux_047:reset, fifo_stage3_to_4:reset_n, fifo_stage3_to_4_in_csr_translator:reset, fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage3_to_4_in_translator:reset, fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:reset, fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage3_to_4_out_translator:reset, fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:reset, fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_046:reset, id_router_047:reset, id_router_053:reset, rsp_xbar_demux_046:reset, rsp_xbar_demux_047:reset, rsp_xbar_demux_053:reset]
	wire          rst_controller_013_reset_out_reset;                                                                 // rst_controller_013:reset_out -> [cmd_xbar_mux_024:reset, fifo_stage4_to_5:reset_n, fifo_stage4_to_5_in_csr_translator:reset, fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage4_to_5_in_translator:reset, fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:reset, fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage4_to_5_out_translator:reset, fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:reset, fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_024:reset, id_router_030:reset, id_router_054:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_054:reset]
	wire          rst_controller_014_reset_out_reset;                                                                 // rst_controller_014:reset_out -> [cmd_xbar_mux_023:reset, fifo_stage5_to_6:reset_n, fifo_stage5_to_6_in_csr_translator:reset, fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage5_to_6_in_translator:reset, fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:reset, fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_stage5_to_6_out_translator:reset, fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:reset, fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_022:reset, id_router_023:reset, id_router_031:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_031:reset]
	wire          rst_controller_015_reset_out_reset;                                                                 // rst_controller_015:reset_out -> [cmd_xbar_mux_001:reset, id_router_001:reset, rsp_xbar_demux_001:reset, sdram_controller:reset_n, sdram_controller_s1_translator:reset, sdram_controller_s1_translator_avalon_universal_slave_0_agent:reset, sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                    // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                          // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                  // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src0_data;                                                                           // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [54:0] cmd_xbar_demux_src0_channel;                                                                        // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                          // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                    // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                          // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                  // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src1_data;                                                                           // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [54:0] cmd_xbar_demux_src1_channel;                                                                        // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                          // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                      // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                              // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src0_data;                                                                       // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [54:0] cmd_xbar_demux_001_src0_channel;                                                                    // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                      // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                      // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                              // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src1_data;                                                                       // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [54:0] cmd_xbar_demux_001_src1_channel;                                                                    // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                      // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                // cmd_xbar_demux_001:src2_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                      // cmd_xbar_demux_001:src2_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                              // cmd_xbar_demux_001:src2_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src2_data;                                                                       // cmd_xbar_demux_001:src2_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_001_src2_channel;                                                                    // cmd_xbar_demux_001:src2_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                // cmd_xbar_demux_001:src3_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                      // cmd_xbar_demux_001:src3_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                              // cmd_xbar_demux_001:src3_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src3_data;                                                                       // cmd_xbar_demux_001:src3_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_001_src3_channel;                                                                    // cmd_xbar_demux_001:src3_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                // cmd_xbar_demux_001:src4_endofpacket -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                      // cmd_xbar_demux_001:src4_valid -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                              // cmd_xbar_demux_001:src4_startofpacket -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src4_data;                                                                       // cmd_xbar_demux_001:src4_data -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_001_src4_channel;                                                                    // cmd_xbar_demux_001:src4_channel -> fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                      // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                              // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src5_data;                                                                       // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [54:0] cmd_xbar_demux_001_src5_channel;                                                                    // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                      // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux_001:src5_ready
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                // cmd_xbar_demux_001:src6_endofpacket -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                      // cmd_xbar_demux_001:src6_valid -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                              // cmd_xbar_demux_001:src6_startofpacket -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src6_data;                                                                       // cmd_xbar_demux_001:src6_data -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_001_src6_channel;                                                                    // cmd_xbar_demux_001:src6_channel -> fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                // cmd_xbar_demux_001:src7_endofpacket -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                      // cmd_xbar_demux_001:src7_valid -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                              // cmd_xbar_demux_001:src7_startofpacket -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src7_data;                                                                       // cmd_xbar_demux_001:src7_data -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_001_src7_channel;                                                                    // cmd_xbar_demux_001:src7_channel -> fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                // cmd_xbar_demux_001:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                      // cmd_xbar_demux_001:src8_valid -> cmd_xbar_mux_008:sink0_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                              // cmd_xbar_demux_001:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src8_data;                                                                       // cmd_xbar_demux_001:src8_data -> cmd_xbar_mux_008:sink0_data
	wire   [54:0] cmd_xbar_demux_001_src8_channel;                                                                    // cmd_xbar_demux_001:src8_channel -> cmd_xbar_mux_008:sink0_channel
	wire          cmd_xbar_demux_001_src8_ready;                                                                      // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux_001:src8_ready
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                // cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                      // cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink0_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                              // cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src9_data;                                                                       // cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink0_data
	wire   [54:0] cmd_xbar_demux_001_src9_channel;                                                                    // cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink0_channel
	wire          cmd_xbar_demux_001_src9_ready;                                                                      // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux_001:src9_ready
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                               // cmd_xbar_demux_001:src10_endofpacket -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                     // cmd_xbar_demux_001:src10_valid -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                             // cmd_xbar_demux_001:src10_startofpacket -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src10_data;                                                                      // cmd_xbar_demux_001:src10_data -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_001_src10_channel;                                                                   // cmd_xbar_demux_001:src10_channel -> fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                               // cmd_xbar_demux_001:src11_endofpacket -> cmd_xbar_mux_011:sink0_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                     // cmd_xbar_demux_001:src11_valid -> cmd_xbar_mux_011:sink0_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                             // cmd_xbar_demux_001:src11_startofpacket -> cmd_xbar_mux_011:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src11_data;                                                                      // cmd_xbar_demux_001:src11_data -> cmd_xbar_mux_011:sink0_data
	wire   [54:0] cmd_xbar_demux_001_src11_channel;                                                                   // cmd_xbar_demux_001:src11_channel -> cmd_xbar_mux_011:sink0_channel
	wire          cmd_xbar_demux_001_src11_ready;                                                                     // cmd_xbar_mux_011:sink0_ready -> cmd_xbar_demux_001:src11_ready
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                               // cmd_xbar_demux_001:src12_endofpacket -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                     // cmd_xbar_demux_001:src12_valid -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                             // cmd_xbar_demux_001:src12_startofpacket -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src12_data;                                                                      // cmd_xbar_demux_001:src12_data -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_001_src12_channel;                                                                   // cmd_xbar_demux_001:src12_channel -> fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                               // cmd_xbar_demux_001:src13_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                     // cmd_xbar_demux_001:src13_valid -> cmd_xbar_mux_013:sink0_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                             // cmd_xbar_demux_001:src13_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src13_data;                                                                      // cmd_xbar_demux_001:src13_data -> cmd_xbar_mux_013:sink0_data
	wire   [54:0] cmd_xbar_demux_001_src13_channel;                                                                   // cmd_xbar_demux_001:src13_channel -> cmd_xbar_mux_013:sink0_channel
	wire          cmd_xbar_demux_001_src13_ready;                                                                     // cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux_001:src13_ready
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                               // cmd_xbar_demux_001:src14_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                     // cmd_xbar_demux_001:src14_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                             // cmd_xbar_demux_001:src14_startofpacket -> width_adapter:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src14_data;                                                                      // cmd_xbar_demux_001:src14_data -> width_adapter:in_data
	wire   [54:0] cmd_xbar_demux_001_src14_channel;                                                                   // cmd_xbar_demux_001:src14_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                               // cmd_xbar_demux_001:src15_endofpacket -> cmd_xbar_mux_015:sink0_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                     // cmd_xbar_demux_001:src15_valid -> cmd_xbar_mux_015:sink0_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                             // cmd_xbar_demux_001:src15_startofpacket -> cmd_xbar_mux_015:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src15_data;                                                                      // cmd_xbar_demux_001:src15_data -> cmd_xbar_mux_015:sink0_data
	wire   [54:0] cmd_xbar_demux_001_src15_channel;                                                                   // cmd_xbar_demux_001:src15_channel -> cmd_xbar_mux_015:sink0_channel
	wire          cmd_xbar_demux_001_src15_ready;                                                                     // cmd_xbar_mux_015:sink0_ready -> cmd_xbar_demux_001:src15_ready
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                               // cmd_xbar_demux_001:src16_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                     // cmd_xbar_demux_001:src16_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                             // cmd_xbar_demux_001:src16_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src16_data;                                                                      // cmd_xbar_demux_001:src16_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_001_src16_channel;                                                                   // cmd_xbar_demux_001:src16_channel -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                      // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_001:sink2_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                              // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src0_data;                                                                       // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_001:sink2_data
	wire   [54:0] cmd_xbar_demux_002_src0_channel;                                                                    // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_001:sink2_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                      // cmd_xbar_mux_001:sink2_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                                // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_015:sink1_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                      // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_015:sink1_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                              // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_015:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src1_data;                                                                       // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_015:sink1_data
	wire   [54:0] cmd_xbar_demux_002_src1_channel;                                                                    // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_015:sink1_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                      // cmd_xbar_mux_015:sink1_ready -> cmd_xbar_demux_002:src1_ready
	wire          cmd_xbar_demux_002_src2_endofpacket;                                                                // cmd_xbar_demux_002:src2_endofpacket -> cmd_xbar_mux_017:sink0_endofpacket
	wire          cmd_xbar_demux_002_src2_valid;                                                                      // cmd_xbar_demux_002:src2_valid -> cmd_xbar_mux_017:sink0_valid
	wire          cmd_xbar_demux_002_src2_startofpacket;                                                              // cmd_xbar_demux_002:src2_startofpacket -> cmd_xbar_mux_017:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src2_data;                                                                       // cmd_xbar_demux_002:src2_data -> cmd_xbar_mux_017:sink0_data
	wire   [54:0] cmd_xbar_demux_002_src2_channel;                                                                    // cmd_xbar_demux_002:src2_channel -> cmd_xbar_mux_017:sink0_channel
	wire          cmd_xbar_demux_002_src2_ready;                                                                      // cmd_xbar_mux_017:sink0_ready -> cmd_xbar_demux_002:src2_ready
	wire          cmd_xbar_demux_002_src3_endofpacket;                                                                // cmd_xbar_demux_002:src3_endofpacket -> cmd_xbar_mux_018:sink0_endofpacket
	wire          cmd_xbar_demux_002_src3_valid;                                                                      // cmd_xbar_demux_002:src3_valid -> cmd_xbar_mux_018:sink0_valid
	wire          cmd_xbar_demux_002_src3_startofpacket;                                                              // cmd_xbar_demux_002:src3_startofpacket -> cmd_xbar_mux_018:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src3_data;                                                                       // cmd_xbar_demux_002:src3_data -> cmd_xbar_mux_018:sink0_data
	wire   [54:0] cmd_xbar_demux_002_src3_channel;                                                                    // cmd_xbar_demux_002:src3_channel -> cmd_xbar_mux_018:sink0_channel
	wire          cmd_xbar_demux_002_src3_ready;                                                                      // cmd_xbar_mux_018:sink0_ready -> cmd_xbar_demux_002:src3_ready
	wire          cmd_xbar_demux_002_src4_endofpacket;                                                                // cmd_xbar_demux_002:src4_endofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src4_valid;                                                                      // cmd_xbar_demux_002:src4_valid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src4_startofpacket;                                                              // cmd_xbar_demux_002:src4_startofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src4_data;                                                                       // cmd_xbar_demux_002:src4_data -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_002_src4_channel;                                                                    // cmd_xbar_demux_002:src4_channel -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src5_endofpacket;                                                                // cmd_xbar_demux_002:src5_endofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src5_valid;                                                                      // cmd_xbar_demux_002:src5_valid -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src5_startofpacket;                                                              // cmd_xbar_demux_002:src5_startofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src5_data;                                                                       // cmd_xbar_demux_002:src5_data -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_002_src5_channel;                                                                    // cmd_xbar_demux_002:src5_channel -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src6_endofpacket;                                                                // cmd_xbar_demux_002:src6_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_002_src6_valid;                                                                      // cmd_xbar_demux_002:src6_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_002_src6_startofpacket;                                                              // cmd_xbar_demux_002:src6_startofpacket -> width_adapter_002:in_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src6_data;                                                                       // cmd_xbar_demux_002:src6_data -> width_adapter_002:in_data
	wire   [54:0] cmd_xbar_demux_002_src6_channel;                                                                    // cmd_xbar_demux_002:src6_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_002_src7_endofpacket;                                                                // cmd_xbar_demux_002:src7_endofpacket -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src7_valid;                                                                      // cmd_xbar_demux_002:src7_valid -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src7_startofpacket;                                                              // cmd_xbar_demux_002:src7_startofpacket -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src7_data;                                                                       // cmd_xbar_demux_002:src7_data -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_002_src7_channel;                                                                    // cmd_xbar_demux_002:src7_channel -> fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src8_endofpacket;                                                                // cmd_xbar_demux_002:src8_endofpacket -> cmd_xbar_mux_023:sink0_endofpacket
	wire          cmd_xbar_demux_002_src8_valid;                                                                      // cmd_xbar_demux_002:src8_valid -> cmd_xbar_mux_023:sink0_valid
	wire          cmd_xbar_demux_002_src8_startofpacket;                                                              // cmd_xbar_demux_002:src8_startofpacket -> cmd_xbar_mux_023:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src8_data;                                                                       // cmd_xbar_demux_002:src8_data -> cmd_xbar_mux_023:sink0_data
	wire   [54:0] cmd_xbar_demux_002_src8_channel;                                                                    // cmd_xbar_demux_002:src8_channel -> cmd_xbar_mux_023:sink0_channel
	wire          cmd_xbar_demux_002_src8_ready;                                                                      // cmd_xbar_mux_023:sink0_ready -> cmd_xbar_demux_002:src8_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_001:sink3_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                      // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_001:sink3_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                              // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_001:sink3_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src0_data;                                                                       // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_001:sink3_data
	wire   [54:0] cmd_xbar_demux_003_src0_channel;                                                                    // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_001:sink3_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                      // cmd_xbar_mux_001:sink3_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                                // cmd_xbar_demux_003:src1_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                      // cmd_xbar_demux_003:src1_valid -> cmd_xbar_mux_013:sink1_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                              // cmd_xbar_demux_003:src1_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src1_data;                                                                       // cmd_xbar_demux_003:src1_data -> cmd_xbar_mux_013:sink1_data
	wire   [54:0] cmd_xbar_demux_003_src1_channel;                                                                    // cmd_xbar_demux_003:src1_channel -> cmd_xbar_mux_013:sink1_channel
	wire          cmd_xbar_demux_003_src1_ready;                                                                      // cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_003:src1_ready
	wire          cmd_xbar_demux_003_src2_endofpacket;                                                                // cmd_xbar_demux_003:src2_endofpacket -> cmd_xbar_mux_023:sink1_endofpacket
	wire          cmd_xbar_demux_003_src2_valid;                                                                      // cmd_xbar_demux_003:src2_valid -> cmd_xbar_mux_023:sink1_valid
	wire          cmd_xbar_demux_003_src2_startofpacket;                                                              // cmd_xbar_demux_003:src2_startofpacket -> cmd_xbar_mux_023:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src2_data;                                                                       // cmd_xbar_demux_003:src2_data -> cmd_xbar_mux_023:sink1_data
	wire   [54:0] cmd_xbar_demux_003_src2_channel;                                                                    // cmd_xbar_demux_003:src2_channel -> cmd_xbar_mux_023:sink1_channel
	wire          cmd_xbar_demux_003_src2_ready;                                                                      // cmd_xbar_mux_023:sink1_ready -> cmd_xbar_demux_003:src2_ready
	wire          cmd_xbar_demux_003_src3_endofpacket;                                                                // cmd_xbar_demux_003:src3_endofpacket -> cmd_xbar_mux_024:sink0_endofpacket
	wire          cmd_xbar_demux_003_src3_valid;                                                                      // cmd_xbar_demux_003:src3_valid -> cmd_xbar_mux_024:sink0_valid
	wire          cmd_xbar_demux_003_src3_startofpacket;                                                              // cmd_xbar_demux_003:src3_startofpacket -> cmd_xbar_mux_024:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src3_data;                                                                       // cmd_xbar_demux_003:src3_data -> cmd_xbar_mux_024:sink0_data
	wire   [54:0] cmd_xbar_demux_003_src3_channel;                                                                    // cmd_xbar_demux_003:src3_channel -> cmd_xbar_mux_024:sink0_channel
	wire          cmd_xbar_demux_003_src3_ready;                                                                      // cmd_xbar_mux_024:sink0_ready -> cmd_xbar_demux_003:src3_ready
	wire          cmd_xbar_demux_003_src4_endofpacket;                                                                // cmd_xbar_demux_003:src4_endofpacket -> cmd_xbar_mux_025:sink0_endofpacket
	wire          cmd_xbar_demux_003_src4_valid;                                                                      // cmd_xbar_demux_003:src4_valid -> cmd_xbar_mux_025:sink0_valid
	wire          cmd_xbar_demux_003_src4_startofpacket;                                                              // cmd_xbar_demux_003:src4_startofpacket -> cmd_xbar_mux_025:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src4_data;                                                                       // cmd_xbar_demux_003:src4_data -> cmd_xbar_mux_025:sink0_data
	wire   [54:0] cmd_xbar_demux_003_src4_channel;                                                                    // cmd_xbar_demux_003:src4_channel -> cmd_xbar_mux_025:sink0_channel
	wire          cmd_xbar_demux_003_src4_ready;                                                                      // cmd_xbar_mux_025:sink0_ready -> cmd_xbar_demux_003:src4_ready
	wire          cmd_xbar_demux_003_src5_endofpacket;                                                                // cmd_xbar_demux_003:src5_endofpacket -> cmd_xbar_mux_026:sink0_endofpacket
	wire          cmd_xbar_demux_003_src5_valid;                                                                      // cmd_xbar_demux_003:src5_valid -> cmd_xbar_mux_026:sink0_valid
	wire          cmd_xbar_demux_003_src5_startofpacket;                                                              // cmd_xbar_demux_003:src5_startofpacket -> cmd_xbar_mux_026:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src5_data;                                                                       // cmd_xbar_demux_003:src5_data -> cmd_xbar_mux_026:sink0_data
	wire   [54:0] cmd_xbar_demux_003_src5_channel;                                                                    // cmd_xbar_demux_003:src5_channel -> cmd_xbar_mux_026:sink0_channel
	wire          cmd_xbar_demux_003_src5_ready;                                                                      // cmd_xbar_mux_026:sink0_ready -> cmd_xbar_demux_003:src5_ready
	wire          cmd_xbar_demux_003_src6_endofpacket;                                                                // cmd_xbar_demux_003:src6_endofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src6_valid;                                                                      // cmd_xbar_demux_003:src6_valid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src6_startofpacket;                                                              // cmd_xbar_demux_003:src6_startofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src6_data;                                                                       // cmd_xbar_demux_003:src6_data -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_003_src6_channel;                                                                    // cmd_xbar_demux_003:src6_channel -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src7_endofpacket;                                                                // cmd_xbar_demux_003:src7_endofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src7_valid;                                                                      // cmd_xbar_demux_003:src7_valid -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src7_startofpacket;                                                              // cmd_xbar_demux_003:src7_startofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src7_data;                                                                       // cmd_xbar_demux_003:src7_data -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_003_src7_channel;                                                                    // cmd_xbar_demux_003:src7_channel -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src8_endofpacket;                                                                // cmd_xbar_demux_003:src8_endofpacket -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src8_valid;                                                                      // cmd_xbar_demux_003:src8_valid -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src8_startofpacket;                                                              // cmd_xbar_demux_003:src8_startofpacket -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src8_data;                                                                       // cmd_xbar_demux_003:src8_data -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_003_src8_channel;                                                                    // cmd_xbar_demux_003:src8_channel -> fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src9_endofpacket;                                                                // cmd_xbar_demux_003:src9_endofpacket -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src9_valid;                                                                      // cmd_xbar_demux_003:src9_valid -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src9_startofpacket;                                                              // cmd_xbar_demux_003:src9_startofpacket -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src9_data;                                                                       // cmd_xbar_demux_003:src9_data -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_003_src9_channel;                                                                    // cmd_xbar_demux_003:src9_channel -> fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src10_endofpacket;                                                               // cmd_xbar_demux_003:src10_endofpacket -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src10_valid;                                                                     // cmd_xbar_demux_003:src10_valid -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src10_startofpacket;                                                             // cmd_xbar_demux_003:src10_startofpacket -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src10_data;                                                                      // cmd_xbar_demux_003:src10_data -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_003_src10_channel;                                                                   // cmd_xbar_demux_003:src10_channel -> fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_001:sink4_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                      // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_001:sink4_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                              // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_001:sink4_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src0_data;                                                                       // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_001:sink4_data
	wire   [54:0] cmd_xbar_demux_004_src0_channel;                                                                    // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_001:sink4_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                      // cmd_xbar_mux_001:sink4_ready -> cmd_xbar_demux_004:src0_ready
	wire          cmd_xbar_demux_004_src1_endofpacket;                                                                // cmd_xbar_demux_004:src1_endofpacket -> cmd_xbar_mux_025:sink1_endofpacket
	wire          cmd_xbar_demux_004_src1_valid;                                                                      // cmd_xbar_demux_004:src1_valid -> cmd_xbar_mux_025:sink1_valid
	wire          cmd_xbar_demux_004_src1_startofpacket;                                                              // cmd_xbar_demux_004:src1_startofpacket -> cmd_xbar_mux_025:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src1_data;                                                                       // cmd_xbar_demux_004:src1_data -> cmd_xbar_mux_025:sink1_data
	wire   [54:0] cmd_xbar_demux_004_src1_channel;                                                                    // cmd_xbar_demux_004:src1_channel -> cmd_xbar_mux_025:sink1_channel
	wire          cmd_xbar_demux_004_src1_ready;                                                                      // cmd_xbar_mux_025:sink1_ready -> cmd_xbar_demux_004:src1_ready
	wire          cmd_xbar_demux_004_src2_endofpacket;                                                                // cmd_xbar_demux_004:src2_endofpacket -> cmd_xbar_mux_026:sink1_endofpacket
	wire          cmd_xbar_demux_004_src2_valid;                                                                      // cmd_xbar_demux_004:src2_valid -> cmd_xbar_mux_026:sink1_valid
	wire          cmd_xbar_demux_004_src2_startofpacket;                                                              // cmd_xbar_demux_004:src2_startofpacket -> cmd_xbar_mux_026:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src2_data;                                                                       // cmd_xbar_demux_004:src2_data -> cmd_xbar_mux_026:sink1_data
	wire   [54:0] cmd_xbar_demux_004_src2_channel;                                                                    // cmd_xbar_demux_004:src2_channel -> cmd_xbar_mux_026:sink1_channel
	wire          cmd_xbar_demux_004_src2_ready;                                                                      // cmd_xbar_mux_026:sink1_ready -> cmd_xbar_demux_004:src2_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_001:sink5_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                      // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_001:sink5_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                              // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_001:sink5_startofpacket
	wire  [106:0] cmd_xbar_demux_005_src0_data;                                                                       // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_001:sink5_data
	wire   [54:0] cmd_xbar_demux_005_src0_channel;                                                                    // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_001:sink5_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                      // cmd_xbar_mux_001:sink5_ready -> cmd_xbar_demux_005:src0_ready
	wire          cmd_xbar_demux_005_src1_endofpacket;                                                                // cmd_xbar_demux_005:src1_endofpacket -> cmd_xbar_mux_032:sink0_endofpacket
	wire          cmd_xbar_demux_005_src1_valid;                                                                      // cmd_xbar_demux_005:src1_valid -> cmd_xbar_mux_032:sink0_valid
	wire          cmd_xbar_demux_005_src1_startofpacket;                                                              // cmd_xbar_demux_005:src1_startofpacket -> cmd_xbar_mux_032:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_005_src1_data;                                                                       // cmd_xbar_demux_005:src1_data -> cmd_xbar_mux_032:sink0_data
	wire   [54:0] cmd_xbar_demux_005_src1_channel;                                                                    // cmd_xbar_demux_005:src1_channel -> cmd_xbar_mux_032:sink0_channel
	wire          cmd_xbar_demux_005_src1_ready;                                                                      // cmd_xbar_mux_032:sink0_ready -> cmd_xbar_demux_005:src1_ready
	wire          cmd_xbar_demux_005_src2_endofpacket;                                                                // cmd_xbar_demux_005:src2_endofpacket -> cmd_xbar_mux_033:sink0_endofpacket
	wire          cmd_xbar_demux_005_src2_valid;                                                                      // cmd_xbar_demux_005:src2_valid -> cmd_xbar_mux_033:sink0_valid
	wire          cmd_xbar_demux_005_src2_startofpacket;                                                              // cmd_xbar_demux_005:src2_startofpacket -> cmd_xbar_mux_033:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_005_src2_data;                                                                       // cmd_xbar_demux_005:src2_data -> cmd_xbar_mux_033:sink0_data
	wire   [54:0] cmd_xbar_demux_005_src2_channel;                                                                    // cmd_xbar_demux_005:src2_channel -> cmd_xbar_mux_033:sink0_channel
	wire          cmd_xbar_demux_005_src2_ready;                                                                      // cmd_xbar_mux_033:sink0_ready -> cmd_xbar_demux_005:src2_ready
	wire          cmd_xbar_demux_006_src0_endofpacket;                                                                // cmd_xbar_demux_006:src0_endofpacket -> cmd_xbar_mux_001:sink6_endofpacket
	wire          cmd_xbar_demux_006_src0_valid;                                                                      // cmd_xbar_demux_006:src0_valid -> cmd_xbar_mux_001:sink6_valid
	wire          cmd_xbar_demux_006_src0_startofpacket;                                                              // cmd_xbar_demux_006:src0_startofpacket -> cmd_xbar_mux_001:sink6_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src0_data;                                                                       // cmd_xbar_demux_006:src0_data -> cmd_xbar_mux_001:sink6_data
	wire   [54:0] cmd_xbar_demux_006_src0_channel;                                                                    // cmd_xbar_demux_006:src0_channel -> cmd_xbar_mux_001:sink6_channel
	wire          cmd_xbar_demux_006_src0_ready;                                                                      // cmd_xbar_mux_001:sink6_ready -> cmd_xbar_demux_006:src0_ready
	wire          cmd_xbar_demux_006_src1_endofpacket;                                                                // cmd_xbar_demux_006:src1_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_006_src1_valid;                                                                      // cmd_xbar_demux_006:src1_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_006_src1_startofpacket;                                                              // cmd_xbar_demux_006:src1_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src1_data;                                                                       // cmd_xbar_demux_006:src1_data -> cmd_xbar_mux_005:sink1_data
	wire   [54:0] cmd_xbar_demux_006_src1_channel;                                                                    // cmd_xbar_demux_006:src1_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_006_src1_ready;                                                                      // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_006:src1_ready
	wire          cmd_xbar_demux_006_src2_endofpacket;                                                                // cmd_xbar_demux_006:src2_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire          cmd_xbar_demux_006_src2_valid;                                                                      // cmd_xbar_demux_006:src2_valid -> cmd_xbar_mux_008:sink1_valid
	wire          cmd_xbar_demux_006_src2_startofpacket;                                                              // cmd_xbar_demux_006:src2_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src2_data;                                                                       // cmd_xbar_demux_006:src2_data -> cmd_xbar_mux_008:sink1_data
	wire   [54:0] cmd_xbar_demux_006_src2_channel;                                                                    // cmd_xbar_demux_006:src2_channel -> cmd_xbar_mux_008:sink1_channel
	wire          cmd_xbar_demux_006_src2_ready;                                                                      // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_006:src2_ready
	wire          cmd_xbar_demux_006_src3_endofpacket;                                                                // cmd_xbar_demux_006:src3_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire          cmd_xbar_demux_006_src3_valid;                                                                      // cmd_xbar_demux_006:src3_valid -> cmd_xbar_mux_009:sink1_valid
	wire          cmd_xbar_demux_006_src3_startofpacket;                                                              // cmd_xbar_demux_006:src3_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src3_data;                                                                       // cmd_xbar_demux_006:src3_data -> cmd_xbar_mux_009:sink1_data
	wire   [54:0] cmd_xbar_demux_006_src3_channel;                                                                    // cmd_xbar_demux_006:src3_channel -> cmd_xbar_mux_009:sink1_channel
	wire          cmd_xbar_demux_006_src3_ready;                                                                      // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_006:src3_ready
	wire          cmd_xbar_demux_006_src4_endofpacket;                                                                // cmd_xbar_demux_006:src4_endofpacket -> cmd_xbar_mux_032:sink1_endofpacket
	wire          cmd_xbar_demux_006_src4_valid;                                                                      // cmd_xbar_demux_006:src4_valid -> cmd_xbar_mux_032:sink1_valid
	wire          cmd_xbar_demux_006_src4_startofpacket;                                                              // cmd_xbar_demux_006:src4_startofpacket -> cmd_xbar_mux_032:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src4_data;                                                                       // cmd_xbar_demux_006:src4_data -> cmd_xbar_mux_032:sink1_data
	wire   [54:0] cmd_xbar_demux_006_src4_channel;                                                                    // cmd_xbar_demux_006:src4_channel -> cmd_xbar_mux_032:sink1_channel
	wire          cmd_xbar_demux_006_src4_ready;                                                                      // cmd_xbar_mux_032:sink1_ready -> cmd_xbar_demux_006:src4_ready
	wire          cmd_xbar_demux_006_src5_endofpacket;                                                                // cmd_xbar_demux_006:src5_endofpacket -> cmd_xbar_mux_033:sink1_endofpacket
	wire          cmd_xbar_demux_006_src5_valid;                                                                      // cmd_xbar_demux_006:src5_valid -> cmd_xbar_mux_033:sink1_valid
	wire          cmd_xbar_demux_006_src5_startofpacket;                                                              // cmd_xbar_demux_006:src5_startofpacket -> cmd_xbar_mux_033:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src5_data;                                                                       // cmd_xbar_demux_006:src5_data -> cmd_xbar_mux_033:sink1_data
	wire   [54:0] cmd_xbar_demux_006_src5_channel;                                                                    // cmd_xbar_demux_006:src5_channel -> cmd_xbar_mux_033:sink1_channel
	wire          cmd_xbar_demux_006_src5_ready;                                                                      // cmd_xbar_mux_033:sink1_ready -> cmd_xbar_demux_006:src5_ready
	wire          cmd_xbar_demux_006_src6_endofpacket;                                                                // cmd_xbar_demux_006:src6_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_006_src6_valid;                                                                      // cmd_xbar_demux_006:src6_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_006_src6_startofpacket;                                                              // cmd_xbar_demux_006:src6_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src6_data;                                                                       // cmd_xbar_demux_006:src6_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_006_src6_channel;                                                                    // cmd_xbar_demux_006:src6_channel -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_006_src7_endofpacket;                                                                // cmd_xbar_demux_006:src7_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_006_src7_valid;                                                                      // cmd_xbar_demux_006:src7_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_006_src7_startofpacket;                                                              // cmd_xbar_demux_006:src7_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src7_data;                                                                       // cmd_xbar_demux_006:src7_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_006_src7_channel;                                                                    // cmd_xbar_demux_006:src7_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_006_src8_endofpacket;                                                                // cmd_xbar_demux_006:src8_endofpacket -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_006_src8_valid;                                                                      // cmd_xbar_demux_006:src8_valid -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_006_src8_startofpacket;                                                              // cmd_xbar_demux_006:src8_startofpacket -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src8_data;                                                                       // cmd_xbar_demux_006:src8_data -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_006_src8_channel;                                                                    // cmd_xbar_demux_006:src8_channel -> fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_006_src9_endofpacket;                                                                // cmd_xbar_demux_006:src9_endofpacket -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_006_src9_valid;                                                                      // cmd_xbar_demux_006:src9_valid -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_006_src9_startofpacket;                                                              // cmd_xbar_demux_006:src9_startofpacket -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src9_data;                                                                       // cmd_xbar_demux_006:src9_data -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_006_src9_channel;                                                                    // cmd_xbar_demux_006:src9_channel -> fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_006_src10_endofpacket;                                                               // cmd_xbar_demux_006:src10_endofpacket -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_006_src10_valid;                                                                     // cmd_xbar_demux_006:src10_valid -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_006_src10_startofpacket;                                                             // cmd_xbar_demux_006:src10_startofpacket -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src10_data;                                                                      // cmd_xbar_demux_006:src10_data -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_006_src10_channel;                                                                   // cmd_xbar_demux_006:src10_channel -> fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_006_src11_endofpacket;                                                               // cmd_xbar_demux_006:src11_endofpacket -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_006_src11_valid;                                                                     // cmd_xbar_demux_006:src11_valid -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_006_src11_startofpacket;                                                             // cmd_xbar_demux_006:src11_startofpacket -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src11_data;                                                                      // cmd_xbar_demux_006:src11_data -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_006_src11_channel;                                                                   // cmd_xbar_demux_006:src11_channel -> fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_006_src12_endofpacket;                                                               // cmd_xbar_demux_006:src12_endofpacket -> cmd_xbar_mux_040:sink0_endofpacket
	wire          cmd_xbar_demux_006_src12_valid;                                                                     // cmd_xbar_demux_006:src12_valid -> cmd_xbar_mux_040:sink0_valid
	wire          cmd_xbar_demux_006_src12_startofpacket;                                                             // cmd_xbar_demux_006:src12_startofpacket -> cmd_xbar_mux_040:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src12_data;                                                                      // cmd_xbar_demux_006:src12_data -> cmd_xbar_mux_040:sink0_data
	wire   [54:0] cmd_xbar_demux_006_src12_channel;                                                                   // cmd_xbar_demux_006:src12_channel -> cmd_xbar_mux_040:sink0_channel
	wire          cmd_xbar_demux_006_src12_ready;                                                                     // cmd_xbar_mux_040:sink0_ready -> cmd_xbar_demux_006:src12_ready
	wire          cmd_xbar_demux_007_src0_endofpacket;                                                                // cmd_xbar_demux_007:src0_endofpacket -> cmd_xbar_mux_001:sink7_endofpacket
	wire          cmd_xbar_demux_007_src0_valid;                                                                      // cmd_xbar_demux_007:src0_valid -> cmd_xbar_mux_001:sink7_valid
	wire          cmd_xbar_demux_007_src0_startofpacket;                                                              // cmd_xbar_demux_007:src0_startofpacket -> cmd_xbar_mux_001:sink7_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src0_data;                                                                       // cmd_xbar_demux_007:src0_data -> cmd_xbar_mux_001:sink7_data
	wire   [54:0] cmd_xbar_demux_007_src0_channel;                                                                    // cmd_xbar_demux_007:src0_channel -> cmd_xbar_mux_001:sink7_channel
	wire          cmd_xbar_demux_007_src0_ready;                                                                      // cmd_xbar_mux_001:sink7_ready -> cmd_xbar_demux_007:src0_ready
	wire          cmd_xbar_demux_007_src1_endofpacket;                                                                // cmd_xbar_demux_007:src1_endofpacket -> cmd_xbar_mux_040:sink1_endofpacket
	wire          cmd_xbar_demux_007_src1_valid;                                                                      // cmd_xbar_demux_007:src1_valid -> cmd_xbar_mux_040:sink1_valid
	wire          cmd_xbar_demux_007_src1_startofpacket;                                                              // cmd_xbar_demux_007:src1_startofpacket -> cmd_xbar_mux_040:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src1_data;                                                                       // cmd_xbar_demux_007:src1_data -> cmd_xbar_mux_040:sink1_data
	wire   [54:0] cmd_xbar_demux_007_src1_channel;                                                                    // cmd_xbar_demux_007:src1_channel -> cmd_xbar_mux_040:sink1_channel
	wire          cmd_xbar_demux_007_src1_ready;                                                                      // cmd_xbar_mux_040:sink1_ready -> cmd_xbar_demux_007:src1_ready
	wire          cmd_xbar_demux_007_src2_endofpacket;                                                                // cmd_xbar_demux_007:src2_endofpacket -> cmd_xbar_mux_041:sink0_endofpacket
	wire          cmd_xbar_demux_007_src2_valid;                                                                      // cmd_xbar_demux_007:src2_valid -> cmd_xbar_mux_041:sink0_valid
	wire          cmd_xbar_demux_007_src2_startofpacket;                                                              // cmd_xbar_demux_007:src2_startofpacket -> cmd_xbar_mux_041:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src2_data;                                                                       // cmd_xbar_demux_007:src2_data -> cmd_xbar_mux_041:sink0_data
	wire   [54:0] cmd_xbar_demux_007_src2_channel;                                                                    // cmd_xbar_demux_007:src2_channel -> cmd_xbar_mux_041:sink0_channel
	wire          cmd_xbar_demux_007_src2_ready;                                                                      // cmd_xbar_mux_041:sink0_ready -> cmd_xbar_demux_007:src2_ready
	wire          cmd_xbar_demux_007_src3_endofpacket;                                                                // cmd_xbar_demux_007:src3_endofpacket -> cmd_xbar_mux_042:sink0_endofpacket
	wire          cmd_xbar_demux_007_src3_valid;                                                                      // cmd_xbar_demux_007:src3_valid -> cmd_xbar_mux_042:sink0_valid
	wire          cmd_xbar_demux_007_src3_startofpacket;                                                              // cmd_xbar_demux_007:src3_startofpacket -> cmd_xbar_mux_042:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src3_data;                                                                       // cmd_xbar_demux_007:src3_data -> cmd_xbar_mux_042:sink0_data
	wire   [54:0] cmd_xbar_demux_007_src3_channel;                                                                    // cmd_xbar_demux_007:src3_channel -> cmd_xbar_mux_042:sink0_channel
	wire          cmd_xbar_demux_007_src3_ready;                                                                      // cmd_xbar_mux_042:sink0_ready -> cmd_xbar_demux_007:src3_ready
	wire          cmd_xbar_demux_007_src4_endofpacket;                                                                // cmd_xbar_demux_007:src4_endofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src4_valid;                                                                      // cmd_xbar_demux_007:src4_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src4_startofpacket;                                                              // cmd_xbar_demux_007:src4_startofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src4_data;                                                                       // cmd_xbar_demux_007:src4_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_007_src4_channel;                                                                    // cmd_xbar_demux_007:src4_channel -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src5_endofpacket;                                                                // cmd_xbar_demux_007:src5_endofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src5_valid;                                                                      // cmd_xbar_demux_007:src5_valid -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src5_startofpacket;                                                              // cmd_xbar_demux_007:src5_startofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src5_data;                                                                       // cmd_xbar_demux_007:src5_data -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_007_src5_channel;                                                                    // cmd_xbar_demux_007:src5_channel -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src6_endofpacket;                                                                // cmd_xbar_demux_007:src6_endofpacket -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src6_valid;                                                                      // cmd_xbar_demux_007:src6_valid -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src6_startofpacket;                                                              // cmd_xbar_demux_007:src6_startofpacket -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src6_data;                                                                       // cmd_xbar_demux_007:src6_data -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_007_src6_channel;                                                                    // cmd_xbar_demux_007:src6_channel -> fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src7_endofpacket;                                                                // cmd_xbar_demux_007:src7_endofpacket -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src7_valid;                                                                      // cmd_xbar_demux_007:src7_valid -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src7_startofpacket;                                                              // cmd_xbar_demux_007:src7_startofpacket -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src7_data;                                                                       // cmd_xbar_demux_007:src7_data -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_007_src7_channel;                                                                    // cmd_xbar_demux_007:src7_channel -> fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src8_endofpacket;                                                                // cmd_xbar_demux_007:src8_endofpacket -> cmd_xbar_mux_047:sink0_endofpacket
	wire          cmd_xbar_demux_007_src8_valid;                                                                      // cmd_xbar_demux_007:src8_valid -> cmd_xbar_mux_047:sink0_valid
	wire          cmd_xbar_demux_007_src8_startofpacket;                                                              // cmd_xbar_demux_007:src8_startofpacket -> cmd_xbar_mux_047:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src8_data;                                                                       // cmd_xbar_demux_007:src8_data -> cmd_xbar_mux_047:sink0_data
	wire   [54:0] cmd_xbar_demux_007_src8_channel;                                                                    // cmd_xbar_demux_007:src8_channel -> cmd_xbar_mux_047:sink0_channel
	wire          cmd_xbar_demux_007_src8_ready;                                                                      // cmd_xbar_mux_047:sink0_ready -> cmd_xbar_demux_007:src8_ready
	wire          cmd_xbar_demux_008_src0_endofpacket;                                                                // cmd_xbar_demux_008:src0_endofpacket -> cmd_xbar_mux_001:sink8_endofpacket
	wire          cmd_xbar_demux_008_src0_valid;                                                                      // cmd_xbar_demux_008:src0_valid -> cmd_xbar_mux_001:sink8_valid
	wire          cmd_xbar_demux_008_src0_startofpacket;                                                              // cmd_xbar_demux_008:src0_startofpacket -> cmd_xbar_mux_001:sink8_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src0_data;                                                                       // cmd_xbar_demux_008:src0_data -> cmd_xbar_mux_001:sink8_data
	wire   [54:0] cmd_xbar_demux_008_src0_channel;                                                                    // cmd_xbar_demux_008:src0_channel -> cmd_xbar_mux_001:sink8_channel
	wire          cmd_xbar_demux_008_src0_ready;                                                                      // cmd_xbar_mux_001:sink8_ready -> cmd_xbar_demux_008:src0_ready
	wire          cmd_xbar_demux_008_src1_endofpacket;                                                                // cmd_xbar_demux_008:src1_endofpacket -> cmd_xbar_mux_011:sink1_endofpacket
	wire          cmd_xbar_demux_008_src1_valid;                                                                      // cmd_xbar_demux_008:src1_valid -> cmd_xbar_mux_011:sink1_valid
	wire          cmd_xbar_demux_008_src1_startofpacket;                                                              // cmd_xbar_demux_008:src1_startofpacket -> cmd_xbar_mux_011:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src1_data;                                                                       // cmd_xbar_demux_008:src1_data -> cmd_xbar_mux_011:sink1_data
	wire   [54:0] cmd_xbar_demux_008_src1_channel;                                                                    // cmd_xbar_demux_008:src1_channel -> cmd_xbar_mux_011:sink1_channel
	wire          cmd_xbar_demux_008_src1_ready;                                                                      // cmd_xbar_mux_011:sink1_ready -> cmd_xbar_demux_008:src1_ready
	wire          cmd_xbar_demux_008_src2_endofpacket;                                                                // cmd_xbar_demux_008:src2_endofpacket -> cmd_xbar_mux_024:sink1_endofpacket
	wire          cmd_xbar_demux_008_src2_valid;                                                                      // cmd_xbar_demux_008:src2_valid -> cmd_xbar_mux_024:sink1_valid
	wire          cmd_xbar_demux_008_src2_startofpacket;                                                              // cmd_xbar_demux_008:src2_startofpacket -> cmd_xbar_mux_024:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src2_data;                                                                       // cmd_xbar_demux_008:src2_data -> cmd_xbar_mux_024:sink1_data
	wire   [54:0] cmd_xbar_demux_008_src2_channel;                                                                    // cmd_xbar_demux_008:src2_channel -> cmd_xbar_mux_024:sink1_channel
	wire          cmd_xbar_demux_008_src2_ready;                                                                      // cmd_xbar_mux_024:sink1_ready -> cmd_xbar_demux_008:src2_ready
	wire          cmd_xbar_demux_008_src3_endofpacket;                                                                // cmd_xbar_demux_008:src3_endofpacket -> cmd_xbar_mux_047:sink1_endofpacket
	wire          cmd_xbar_demux_008_src3_valid;                                                                      // cmd_xbar_demux_008:src3_valid -> cmd_xbar_mux_047:sink1_valid
	wire          cmd_xbar_demux_008_src3_startofpacket;                                                              // cmd_xbar_demux_008:src3_startofpacket -> cmd_xbar_mux_047:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src3_data;                                                                       // cmd_xbar_demux_008:src3_data -> cmd_xbar_mux_047:sink1_data
	wire   [54:0] cmd_xbar_demux_008_src3_channel;                                                                    // cmd_xbar_demux_008:src3_channel -> cmd_xbar_mux_047:sink1_channel
	wire          cmd_xbar_demux_008_src3_ready;                                                                      // cmd_xbar_mux_047:sink1_ready -> cmd_xbar_demux_008:src3_ready
	wire          cmd_xbar_demux_008_src4_endofpacket;                                                                // cmd_xbar_demux_008:src4_endofpacket -> cmd_xbar_mux_048:sink0_endofpacket
	wire          cmd_xbar_demux_008_src4_valid;                                                                      // cmd_xbar_demux_008:src4_valid -> cmd_xbar_mux_048:sink0_valid
	wire          cmd_xbar_demux_008_src4_startofpacket;                                                              // cmd_xbar_demux_008:src4_startofpacket -> cmd_xbar_mux_048:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src4_data;                                                                       // cmd_xbar_demux_008:src4_data -> cmd_xbar_mux_048:sink0_data
	wire   [54:0] cmd_xbar_demux_008_src4_channel;                                                                    // cmd_xbar_demux_008:src4_channel -> cmd_xbar_mux_048:sink0_channel
	wire          cmd_xbar_demux_008_src4_ready;                                                                      // cmd_xbar_mux_048:sink0_ready -> cmd_xbar_demux_008:src4_ready
	wire          cmd_xbar_demux_008_src5_endofpacket;                                                                // cmd_xbar_demux_008:src5_endofpacket -> cmd_xbar_mux_049:sink0_endofpacket
	wire          cmd_xbar_demux_008_src5_valid;                                                                      // cmd_xbar_demux_008:src5_valid -> cmd_xbar_mux_049:sink0_valid
	wire          cmd_xbar_demux_008_src5_startofpacket;                                                              // cmd_xbar_demux_008:src5_startofpacket -> cmd_xbar_mux_049:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src5_data;                                                                       // cmd_xbar_demux_008:src5_data -> cmd_xbar_mux_049:sink0_data
	wire   [54:0] cmd_xbar_demux_008_src5_channel;                                                                    // cmd_xbar_demux_008:src5_channel -> cmd_xbar_mux_049:sink0_channel
	wire          cmd_xbar_demux_008_src5_ready;                                                                      // cmd_xbar_mux_049:sink0_ready -> cmd_xbar_demux_008:src5_ready
	wire          cmd_xbar_demux_008_src6_endofpacket;                                                                // cmd_xbar_demux_008:src6_endofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src6_valid;                                                                      // cmd_xbar_demux_008:src6_valid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src6_startofpacket;                                                              // cmd_xbar_demux_008:src6_startofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src6_data;                                                                       // cmd_xbar_demux_008:src6_data -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_008_src6_channel;                                                                    // cmd_xbar_demux_008:src6_channel -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src7_endofpacket;                                                                // cmd_xbar_demux_008:src7_endofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src7_valid;                                                                      // cmd_xbar_demux_008:src7_valid -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src7_startofpacket;                                                              // cmd_xbar_demux_008:src7_startofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src7_data;                                                                       // cmd_xbar_demux_008:src7_data -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_008_src7_channel;                                                                    // cmd_xbar_demux_008:src7_channel -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src8_endofpacket;                                                                // cmd_xbar_demux_008:src8_endofpacket -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src8_valid;                                                                      // cmd_xbar_demux_008:src8_valid -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src8_startofpacket;                                                              // cmd_xbar_demux_008:src8_startofpacket -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src8_data;                                                                       // cmd_xbar_demux_008:src8_data -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_008_src8_channel;                                                                    // cmd_xbar_demux_008:src8_channel -> fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src9_endofpacket;                                                                // cmd_xbar_demux_008:src9_endofpacket -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src9_valid;                                                                      // cmd_xbar_demux_008:src9_valid -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src9_startofpacket;                                                              // cmd_xbar_demux_008:src9_startofpacket -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src9_data;                                                                       // cmd_xbar_demux_008:src9_data -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_008_src9_channel;                                                                    // cmd_xbar_demux_008:src9_channel -> fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src10_endofpacket;                                                               // cmd_xbar_demux_008:src10_endofpacket -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src10_valid;                                                                     // cmd_xbar_demux_008:src10_valid -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src10_startofpacket;                                                             // cmd_xbar_demux_008:src10_startofpacket -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src10_data;                                                                      // cmd_xbar_demux_008:src10_data -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_demux_008_src10_channel;                                                                   // cmd_xbar_demux_008:src10_channel -> fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_009_src0_endofpacket;                                                                // cmd_xbar_demux_009:src0_endofpacket -> cmd_xbar_mux_001:sink9_endofpacket
	wire          cmd_xbar_demux_009_src0_valid;                                                                      // cmd_xbar_demux_009:src0_valid -> cmd_xbar_mux_001:sink9_valid
	wire          cmd_xbar_demux_009_src0_startofpacket;                                                              // cmd_xbar_demux_009:src0_startofpacket -> cmd_xbar_mux_001:sink9_startofpacket
	wire  [106:0] cmd_xbar_demux_009_src0_data;                                                                       // cmd_xbar_demux_009:src0_data -> cmd_xbar_mux_001:sink9_data
	wire   [54:0] cmd_xbar_demux_009_src0_channel;                                                                    // cmd_xbar_demux_009:src0_channel -> cmd_xbar_mux_001:sink9_channel
	wire          cmd_xbar_demux_009_src0_ready;                                                                      // cmd_xbar_mux_001:sink9_ready -> cmd_xbar_demux_009:src0_ready
	wire          cmd_xbar_demux_009_src1_endofpacket;                                                                // cmd_xbar_demux_009:src1_endofpacket -> cmd_xbar_mux_048:sink1_endofpacket
	wire          cmd_xbar_demux_009_src1_valid;                                                                      // cmd_xbar_demux_009:src1_valid -> cmd_xbar_mux_048:sink1_valid
	wire          cmd_xbar_demux_009_src1_startofpacket;                                                              // cmd_xbar_demux_009:src1_startofpacket -> cmd_xbar_mux_048:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_009_src1_data;                                                                       // cmd_xbar_demux_009:src1_data -> cmd_xbar_mux_048:sink1_data
	wire   [54:0] cmd_xbar_demux_009_src1_channel;                                                                    // cmd_xbar_demux_009:src1_channel -> cmd_xbar_mux_048:sink1_channel
	wire          cmd_xbar_demux_009_src1_ready;                                                                      // cmd_xbar_mux_048:sink1_ready -> cmd_xbar_demux_009:src1_ready
	wire          cmd_xbar_demux_009_src2_endofpacket;                                                                // cmd_xbar_demux_009:src2_endofpacket -> cmd_xbar_mux_049:sink1_endofpacket
	wire          cmd_xbar_demux_009_src2_valid;                                                                      // cmd_xbar_demux_009:src2_valid -> cmd_xbar_mux_049:sink1_valid
	wire          cmd_xbar_demux_009_src2_startofpacket;                                                              // cmd_xbar_demux_009:src2_startofpacket -> cmd_xbar_mux_049:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_009_src2_data;                                                                       // cmd_xbar_demux_009:src2_data -> cmd_xbar_mux_049:sink1_data
	wire   [54:0] cmd_xbar_demux_009_src2_channel;                                                                    // cmd_xbar_demux_009:src2_channel -> cmd_xbar_mux_049:sink1_channel
	wire          cmd_xbar_demux_009_src2_ready;                                                                      // cmd_xbar_mux_049:sink1_ready -> cmd_xbar_demux_009:src2_ready
	wire          cmd_xbar_demux_010_src0_endofpacket;                                                                // cmd_xbar_demux_010:src0_endofpacket -> cmd_xbar_mux_001:sink10_endofpacket
	wire          cmd_xbar_demux_010_src0_valid;                                                                      // cmd_xbar_demux_010:src0_valid -> cmd_xbar_mux_001:sink10_valid
	wire          cmd_xbar_demux_010_src0_startofpacket;                                                              // cmd_xbar_demux_010:src0_startofpacket -> cmd_xbar_mux_001:sink10_startofpacket
	wire  [106:0] cmd_xbar_demux_010_src0_data;                                                                       // cmd_xbar_demux_010:src0_data -> cmd_xbar_mux_001:sink10_data
	wire   [54:0] cmd_xbar_demux_010_src0_channel;                                                                    // cmd_xbar_demux_010:src0_channel -> cmd_xbar_mux_001:sink10_channel
	wire          cmd_xbar_demux_010_src0_ready;                                                                      // cmd_xbar_mux_001:sink10_ready -> cmd_xbar_demux_010:src0_ready
	wire          cmd_xbar_demux_010_src1_endofpacket;                                                                // cmd_xbar_demux_010:src1_endofpacket -> cmd_xbar_mux_041:sink1_endofpacket
	wire          cmd_xbar_demux_010_src1_valid;                                                                      // cmd_xbar_demux_010:src1_valid -> cmd_xbar_mux_041:sink1_valid
	wire          cmd_xbar_demux_010_src1_startofpacket;                                                              // cmd_xbar_demux_010:src1_startofpacket -> cmd_xbar_mux_041:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_010_src1_data;                                                                       // cmd_xbar_demux_010:src1_data -> cmd_xbar_mux_041:sink1_data
	wire   [54:0] cmd_xbar_demux_010_src1_channel;                                                                    // cmd_xbar_demux_010:src1_channel -> cmd_xbar_mux_041:sink1_channel
	wire          cmd_xbar_demux_010_src1_ready;                                                                      // cmd_xbar_mux_041:sink1_ready -> cmd_xbar_demux_010:src1_ready
	wire          cmd_xbar_demux_010_src2_endofpacket;                                                                // cmd_xbar_demux_010:src2_endofpacket -> cmd_xbar_mux_042:sink1_endofpacket
	wire          cmd_xbar_demux_010_src2_valid;                                                                      // cmd_xbar_demux_010:src2_valid -> cmd_xbar_mux_042:sink1_valid
	wire          cmd_xbar_demux_010_src2_startofpacket;                                                              // cmd_xbar_demux_010:src2_startofpacket -> cmd_xbar_mux_042:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_010_src2_data;                                                                       // cmd_xbar_demux_010:src2_data -> cmd_xbar_mux_042:sink1_data
	wire   [54:0] cmd_xbar_demux_010_src2_channel;                                                                    // cmd_xbar_demux_010:src2_channel -> cmd_xbar_mux_042:sink1_channel
	wire          cmd_xbar_demux_010_src2_ready;                                                                      // cmd_xbar_mux_042:sink1_ready -> cmd_xbar_demux_010:src2_ready
	wire          cmd_xbar_demux_011_src0_endofpacket;                                                                // cmd_xbar_demux_011:src0_endofpacket -> cmd_xbar_mux_001:sink11_endofpacket
	wire          cmd_xbar_demux_011_src0_valid;                                                                      // cmd_xbar_demux_011:src0_valid -> cmd_xbar_mux_001:sink11_valid
	wire          cmd_xbar_demux_011_src0_startofpacket;                                                              // cmd_xbar_demux_011:src0_startofpacket -> cmd_xbar_mux_001:sink11_startofpacket
	wire  [106:0] cmd_xbar_demux_011_src0_data;                                                                       // cmd_xbar_demux_011:src0_data -> cmd_xbar_mux_001:sink11_data
	wire   [54:0] cmd_xbar_demux_011_src0_channel;                                                                    // cmd_xbar_demux_011:src0_channel -> cmd_xbar_mux_001:sink11_channel
	wire          cmd_xbar_demux_011_src0_ready;                                                                      // cmd_xbar_mux_001:sink11_ready -> cmd_xbar_demux_011:src0_ready
	wire          cmd_xbar_demux_011_src1_endofpacket;                                                                // cmd_xbar_demux_011:src1_endofpacket -> cmd_xbar_mux_017:sink1_endofpacket
	wire          cmd_xbar_demux_011_src1_valid;                                                                      // cmd_xbar_demux_011:src1_valid -> cmd_xbar_mux_017:sink1_valid
	wire          cmd_xbar_demux_011_src1_startofpacket;                                                              // cmd_xbar_demux_011:src1_startofpacket -> cmd_xbar_mux_017:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_011_src1_data;                                                                       // cmd_xbar_demux_011:src1_data -> cmd_xbar_mux_017:sink1_data
	wire   [54:0] cmd_xbar_demux_011_src1_channel;                                                                    // cmd_xbar_demux_011:src1_channel -> cmd_xbar_mux_017:sink1_channel
	wire          cmd_xbar_demux_011_src1_ready;                                                                      // cmd_xbar_mux_017:sink1_ready -> cmd_xbar_demux_011:src1_ready
	wire          cmd_xbar_demux_011_src2_endofpacket;                                                                // cmd_xbar_demux_011:src2_endofpacket -> cmd_xbar_mux_018:sink1_endofpacket
	wire          cmd_xbar_demux_011_src2_valid;                                                                      // cmd_xbar_demux_011:src2_valid -> cmd_xbar_mux_018:sink1_valid
	wire          cmd_xbar_demux_011_src2_startofpacket;                                                              // cmd_xbar_demux_011:src2_startofpacket -> cmd_xbar_mux_018:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_011_src2_data;                                                                       // cmd_xbar_demux_011:src2_data -> cmd_xbar_mux_018:sink1_data
	wire   [54:0] cmd_xbar_demux_011_src2_channel;                                                                    // cmd_xbar_demux_011:src2_channel -> cmd_xbar_mux_018:sink1_channel
	wire          cmd_xbar_demux_011_src2_ready;                                                                      // cmd_xbar_mux_018:sink1_ready -> cmd_xbar_demux_011:src2_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                    // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                          // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                  // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src0_data;                                                                           // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [54:0] rsp_xbar_demux_src0_channel;                                                                        // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                          // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                    // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                          // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                  // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src1_data;                                                                           // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [54:0] rsp_xbar_demux_src1_channel;                                                                        // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                          // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                      // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                              // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src0_data;                                                                       // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [54:0] rsp_xbar_demux_001_src0_channel;                                                                    // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                      // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                      // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                              // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src1_data;                                                                       // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [54:0] rsp_xbar_demux_001_src1_channel;                                                                    // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                      // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                                // rsp_xbar_demux_001:src2_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                      // rsp_xbar_demux_001:src2_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                              // rsp_xbar_demux_001:src2_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src2_data;                                                                       // rsp_xbar_demux_001:src2_data -> rsp_xbar_mux_002:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src2_channel;                                                                    // rsp_xbar_demux_001:src2_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_001_src2_ready;                                                                      // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_001:src2_ready
	wire          rsp_xbar_demux_001_src3_endofpacket;                                                                // rsp_xbar_demux_001:src3_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          rsp_xbar_demux_001_src3_valid;                                                                      // rsp_xbar_demux_001:src3_valid -> rsp_xbar_mux_003:sink0_valid
	wire          rsp_xbar_demux_001_src3_startofpacket;                                                              // rsp_xbar_demux_001:src3_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src3_data;                                                                       // rsp_xbar_demux_001:src3_data -> rsp_xbar_mux_003:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src3_channel;                                                                    // rsp_xbar_demux_001:src3_channel -> rsp_xbar_mux_003:sink0_channel
	wire          rsp_xbar_demux_001_src3_ready;                                                                      // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_001:src3_ready
	wire          rsp_xbar_demux_001_src4_endofpacket;                                                                // rsp_xbar_demux_001:src4_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	wire          rsp_xbar_demux_001_src4_valid;                                                                      // rsp_xbar_demux_001:src4_valid -> rsp_xbar_mux_004:sink0_valid
	wire          rsp_xbar_demux_001_src4_startofpacket;                                                              // rsp_xbar_demux_001:src4_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src4_data;                                                                       // rsp_xbar_demux_001:src4_data -> rsp_xbar_mux_004:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src4_channel;                                                                    // rsp_xbar_demux_001:src4_channel -> rsp_xbar_mux_004:sink0_channel
	wire          rsp_xbar_demux_001_src4_ready;                                                                      // rsp_xbar_mux_004:sink0_ready -> rsp_xbar_demux_001:src4_ready
	wire          rsp_xbar_demux_001_src5_endofpacket;                                                                // rsp_xbar_demux_001:src5_endofpacket -> rsp_xbar_mux_005:sink0_endofpacket
	wire          rsp_xbar_demux_001_src5_valid;                                                                      // rsp_xbar_demux_001:src5_valid -> rsp_xbar_mux_005:sink0_valid
	wire          rsp_xbar_demux_001_src5_startofpacket;                                                              // rsp_xbar_demux_001:src5_startofpacket -> rsp_xbar_mux_005:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src5_data;                                                                       // rsp_xbar_demux_001:src5_data -> rsp_xbar_mux_005:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src5_channel;                                                                    // rsp_xbar_demux_001:src5_channel -> rsp_xbar_mux_005:sink0_channel
	wire          rsp_xbar_demux_001_src5_ready;                                                                      // rsp_xbar_mux_005:sink0_ready -> rsp_xbar_demux_001:src5_ready
	wire          rsp_xbar_demux_001_src6_endofpacket;                                                                // rsp_xbar_demux_001:src6_endofpacket -> rsp_xbar_mux_006:sink0_endofpacket
	wire          rsp_xbar_demux_001_src6_valid;                                                                      // rsp_xbar_demux_001:src6_valid -> rsp_xbar_mux_006:sink0_valid
	wire          rsp_xbar_demux_001_src6_startofpacket;                                                              // rsp_xbar_demux_001:src6_startofpacket -> rsp_xbar_mux_006:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src6_data;                                                                       // rsp_xbar_demux_001:src6_data -> rsp_xbar_mux_006:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src6_channel;                                                                    // rsp_xbar_demux_001:src6_channel -> rsp_xbar_mux_006:sink0_channel
	wire          rsp_xbar_demux_001_src6_ready;                                                                      // rsp_xbar_mux_006:sink0_ready -> rsp_xbar_demux_001:src6_ready
	wire          rsp_xbar_demux_001_src7_endofpacket;                                                                // rsp_xbar_demux_001:src7_endofpacket -> rsp_xbar_mux_007:sink0_endofpacket
	wire          rsp_xbar_demux_001_src7_valid;                                                                      // rsp_xbar_demux_001:src7_valid -> rsp_xbar_mux_007:sink0_valid
	wire          rsp_xbar_demux_001_src7_startofpacket;                                                              // rsp_xbar_demux_001:src7_startofpacket -> rsp_xbar_mux_007:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src7_data;                                                                       // rsp_xbar_demux_001:src7_data -> rsp_xbar_mux_007:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src7_channel;                                                                    // rsp_xbar_demux_001:src7_channel -> rsp_xbar_mux_007:sink0_channel
	wire          rsp_xbar_demux_001_src7_ready;                                                                      // rsp_xbar_mux_007:sink0_ready -> rsp_xbar_demux_001:src7_ready
	wire          rsp_xbar_demux_001_src8_endofpacket;                                                                // rsp_xbar_demux_001:src8_endofpacket -> rsp_xbar_mux_008:sink0_endofpacket
	wire          rsp_xbar_demux_001_src8_valid;                                                                      // rsp_xbar_demux_001:src8_valid -> rsp_xbar_mux_008:sink0_valid
	wire          rsp_xbar_demux_001_src8_startofpacket;                                                              // rsp_xbar_demux_001:src8_startofpacket -> rsp_xbar_mux_008:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src8_data;                                                                       // rsp_xbar_demux_001:src8_data -> rsp_xbar_mux_008:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src8_channel;                                                                    // rsp_xbar_demux_001:src8_channel -> rsp_xbar_mux_008:sink0_channel
	wire          rsp_xbar_demux_001_src8_ready;                                                                      // rsp_xbar_mux_008:sink0_ready -> rsp_xbar_demux_001:src8_ready
	wire          rsp_xbar_demux_001_src9_endofpacket;                                                                // rsp_xbar_demux_001:src9_endofpacket -> rsp_xbar_mux_009:sink0_endofpacket
	wire          rsp_xbar_demux_001_src9_valid;                                                                      // rsp_xbar_demux_001:src9_valid -> rsp_xbar_mux_009:sink0_valid
	wire          rsp_xbar_demux_001_src9_startofpacket;                                                              // rsp_xbar_demux_001:src9_startofpacket -> rsp_xbar_mux_009:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src9_data;                                                                       // rsp_xbar_demux_001:src9_data -> rsp_xbar_mux_009:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src9_channel;                                                                    // rsp_xbar_demux_001:src9_channel -> rsp_xbar_mux_009:sink0_channel
	wire          rsp_xbar_demux_001_src9_ready;                                                                      // rsp_xbar_mux_009:sink0_ready -> rsp_xbar_demux_001:src9_ready
	wire          rsp_xbar_demux_001_src10_endofpacket;                                                               // rsp_xbar_demux_001:src10_endofpacket -> rsp_xbar_mux_010:sink0_endofpacket
	wire          rsp_xbar_demux_001_src10_valid;                                                                     // rsp_xbar_demux_001:src10_valid -> rsp_xbar_mux_010:sink0_valid
	wire          rsp_xbar_demux_001_src10_startofpacket;                                                             // rsp_xbar_demux_001:src10_startofpacket -> rsp_xbar_mux_010:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src10_data;                                                                      // rsp_xbar_demux_001:src10_data -> rsp_xbar_mux_010:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src10_channel;                                                                   // rsp_xbar_demux_001:src10_channel -> rsp_xbar_mux_010:sink0_channel
	wire          rsp_xbar_demux_001_src10_ready;                                                                     // rsp_xbar_mux_010:sink0_ready -> rsp_xbar_demux_001:src10_ready
	wire          rsp_xbar_demux_001_src11_endofpacket;                                                               // rsp_xbar_demux_001:src11_endofpacket -> rsp_xbar_mux_011:sink0_endofpacket
	wire          rsp_xbar_demux_001_src11_valid;                                                                     // rsp_xbar_demux_001:src11_valid -> rsp_xbar_mux_011:sink0_valid
	wire          rsp_xbar_demux_001_src11_startofpacket;                                                             // rsp_xbar_demux_001:src11_startofpacket -> rsp_xbar_mux_011:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src11_data;                                                                      // rsp_xbar_demux_001:src11_data -> rsp_xbar_mux_011:sink0_data
	wire   [54:0] rsp_xbar_demux_001_src11_channel;                                                                   // rsp_xbar_demux_001:src11_channel -> rsp_xbar_mux_011:sink0_channel
	wire          rsp_xbar_demux_001_src11_ready;                                                                     // rsp_xbar_mux_011:sink0_ready -> rsp_xbar_demux_001:src11_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                      // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                              // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src0_data;                                                                       // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire   [54:0] rsp_xbar_demux_002_src0_channel;                                                                    // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                      // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                      // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                              // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src0_data;                                                                       // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [54:0] rsp_xbar_demux_003_src0_channel;                                                                    // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                      // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                      // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                              // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src0_data;                                                                       // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [54:0] rsp_xbar_demux_004_src0_channel;                                                                    // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                      // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                      // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                              // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_005_src0_data;                                                                       // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [54:0] rsp_xbar_demux_005_src0_channel;                                                                    // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                      // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_006:sink1_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                      // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_006:sink1_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                              // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_006:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_005_src1_data;                                                                       // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_006:sink1_data
	wire   [54:0] rsp_xbar_demux_005_src1_channel;                                                                    // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_006:sink1_channel
	wire          rsp_xbar_demux_005_src1_ready;                                                                      // rsp_xbar_mux_006:sink1_ready -> rsp_xbar_demux_005:src1_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                      // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                              // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_006_src0_data;                                                                       // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [54:0] rsp_xbar_demux_006_src0_channel;                                                                    // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                      // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                      // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                              // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_007_src0_data;                                                                       // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [54:0] rsp_xbar_demux_007_src0_channel;                                                                    // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                      // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                      // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                              // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_008_src0_data;                                                                       // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [54:0] rsp_xbar_demux_008_src0_channel;                                                                    // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                      // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_008_src1_endofpacket;                                                                // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_006:sink2_endofpacket
	wire          rsp_xbar_demux_008_src1_valid;                                                                      // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_006:sink2_valid
	wire          rsp_xbar_demux_008_src1_startofpacket;                                                              // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_006:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_008_src1_data;                                                                       // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_006:sink2_data
	wire   [54:0] rsp_xbar_demux_008_src1_channel;                                                                    // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_006:sink2_channel
	wire          rsp_xbar_demux_008_src1_ready;                                                                      // rsp_xbar_mux_006:sink2_ready -> rsp_xbar_demux_008:src1_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                      // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                              // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src0_data;                                                                       // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [54:0] rsp_xbar_demux_009_src0_channel;                                                                    // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                      // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_009_src1_endofpacket;                                                                // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_006:sink3_endofpacket
	wire          rsp_xbar_demux_009_src1_valid;                                                                      // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_006:sink3_valid
	wire          rsp_xbar_demux_009_src1_startofpacket;                                                              // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_006:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src1_data;                                                                       // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_006:sink3_data
	wire   [54:0] rsp_xbar_demux_009_src1_channel;                                                                    // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_006:sink3_channel
	wire          rsp_xbar_demux_009_src1_ready;                                                                      // rsp_xbar_mux_006:sink3_ready -> rsp_xbar_demux_009:src1_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                      // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                              // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [106:0] rsp_xbar_demux_010_src0_data;                                                                       // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [54:0] rsp_xbar_demux_010_src0_channel;                                                                    // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                      // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                      // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                              // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [106:0] rsp_xbar_demux_011_src0_data;                                                                       // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [54:0] rsp_xbar_demux_011_src0_channel;                                                                    // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                      // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_011_src1_endofpacket;                                                                // rsp_xbar_demux_011:src1_endofpacket -> rsp_xbar_mux_008:sink1_endofpacket
	wire          rsp_xbar_demux_011_src1_valid;                                                                      // rsp_xbar_demux_011:src1_valid -> rsp_xbar_mux_008:sink1_valid
	wire          rsp_xbar_demux_011_src1_startofpacket;                                                              // rsp_xbar_demux_011:src1_startofpacket -> rsp_xbar_mux_008:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_011_src1_data;                                                                       // rsp_xbar_demux_011:src1_data -> rsp_xbar_mux_008:sink1_data
	wire   [54:0] rsp_xbar_demux_011_src1_channel;                                                                    // rsp_xbar_demux_011:src1_channel -> rsp_xbar_mux_008:sink1_channel
	wire          rsp_xbar_demux_011_src1_ready;                                                                      // rsp_xbar_mux_008:sink1_ready -> rsp_xbar_demux_011:src1_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                      // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                              // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [106:0] rsp_xbar_demux_012_src0_data;                                                                       // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [54:0] rsp_xbar_demux_012_src0_channel;                                                                    // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                      // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                      // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                              // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src0_data;                                                                       // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [54:0] rsp_xbar_demux_013_src0_channel;                                                                    // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                      // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_013_src1_endofpacket;                                                                // rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          rsp_xbar_demux_013_src1_valid;                                                                      // rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_003:sink1_valid
	wire          rsp_xbar_demux_013_src1_startofpacket;                                                              // rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src1_data;                                                                       // rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_003:sink1_data
	wire   [54:0] rsp_xbar_demux_013_src1_channel;                                                                    // rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_003:sink1_channel
	wire          rsp_xbar_demux_013_src1_ready;                                                                      // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_013:src1_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                      // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                              // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [106:0] rsp_xbar_demux_014_src0_data;                                                                       // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire   [54:0] rsp_xbar_demux_014_src0_channel;                                                                    // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                      // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                      // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                              // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [106:0] rsp_xbar_demux_015_src0_data;                                                                       // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [54:0] rsp_xbar_demux_015_src0_channel;                                                                    // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                      // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_015_src1_endofpacket;                                                                // rsp_xbar_demux_015:src1_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          rsp_xbar_demux_015_src1_valid;                                                                      // rsp_xbar_demux_015:src1_valid -> rsp_xbar_mux_002:sink1_valid
	wire          rsp_xbar_demux_015_src1_startofpacket;                                                              // rsp_xbar_demux_015:src1_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_015_src1_data;                                                                       // rsp_xbar_demux_015:src1_data -> rsp_xbar_mux_002:sink1_data
	wire   [54:0] rsp_xbar_demux_015_src1_channel;                                                                    // rsp_xbar_demux_015:src1_channel -> rsp_xbar_mux_002:sink1_channel
	wire          rsp_xbar_demux_015_src1_ready;                                                                      // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_015:src1_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                      // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                              // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [106:0] rsp_xbar_demux_016_src0_data;                                                                       // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire   [54:0] rsp_xbar_demux_016_src0_channel;                                                                    // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                      // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                      // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_002:sink2_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                              // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_017_src0_data;                                                                       // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_002:sink2_data
	wire   [54:0] rsp_xbar_demux_017_src0_channel;                                                                    // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_002:sink2_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                      // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_017_src1_endofpacket;                                                                // rsp_xbar_demux_017:src1_endofpacket -> rsp_xbar_mux_011:sink1_endofpacket
	wire          rsp_xbar_demux_017_src1_valid;                                                                      // rsp_xbar_demux_017:src1_valid -> rsp_xbar_mux_011:sink1_valid
	wire          rsp_xbar_demux_017_src1_startofpacket;                                                              // rsp_xbar_demux_017:src1_startofpacket -> rsp_xbar_mux_011:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_017_src1_data;                                                                       // rsp_xbar_demux_017:src1_data -> rsp_xbar_mux_011:sink1_data
	wire   [54:0] rsp_xbar_demux_017_src1_channel;                                                                    // rsp_xbar_demux_017:src1_channel -> rsp_xbar_mux_011:sink1_channel
	wire          rsp_xbar_demux_017_src1_ready;                                                                      // rsp_xbar_mux_011:sink1_ready -> rsp_xbar_demux_017:src1_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                      // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_002:sink3_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                              // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_018_src0_data;                                                                       // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_002:sink3_data
	wire   [54:0] rsp_xbar_demux_018_src0_channel;                                                                    // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_002:sink3_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                      // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_018_src1_endofpacket;                                                                // rsp_xbar_demux_018:src1_endofpacket -> rsp_xbar_mux_011:sink2_endofpacket
	wire          rsp_xbar_demux_018_src1_valid;                                                                      // rsp_xbar_demux_018:src1_valid -> rsp_xbar_mux_011:sink2_valid
	wire          rsp_xbar_demux_018_src1_startofpacket;                                                              // rsp_xbar_demux_018:src1_startofpacket -> rsp_xbar_mux_011:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_018_src1_data;                                                                       // rsp_xbar_demux_018:src1_data -> rsp_xbar_mux_011:sink2_data
	wire   [54:0] rsp_xbar_demux_018_src1_channel;                                                                    // rsp_xbar_demux_018:src1_channel -> rsp_xbar_mux_011:sink2_channel
	wire          rsp_xbar_demux_018_src1_ready;                                                                      // rsp_xbar_mux_011:sink2_ready -> rsp_xbar_demux_018:src1_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                      // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_002:sink4_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                              // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_019_src0_data;                                                                       // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_002:sink4_data
	wire   [54:0] rsp_xbar_demux_019_src0_channel;                                                                    // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_002:sink4_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                      // rsp_xbar_mux_002:sink4_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                                // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_002:sink5_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                      // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_002:sink5_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                              // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_002:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_020_src0_data;                                                                       // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_002:sink5_data
	wire   [54:0] rsp_xbar_demux_020_src0_channel;                                                                    // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_002:sink5_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                      // rsp_xbar_mux_002:sink5_ready -> rsp_xbar_demux_020:src0_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                                // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_002:sink6_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                      // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_002:sink6_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                              // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_002:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_021_src0_data;                                                                       // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_002:sink6_data
	wire   [54:0] rsp_xbar_demux_021_src0_channel;                                                                    // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_002:sink6_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                      // rsp_xbar_mux_002:sink6_ready -> rsp_xbar_demux_021:src0_ready
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                                // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_002:sink7_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                      // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_002:sink7_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                              // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_002:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_022_src0_data;                                                                       // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_002:sink7_data
	wire   [54:0] rsp_xbar_demux_022_src0_channel;                                                                    // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_002:sink7_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                      // rsp_xbar_mux_002:sink7_ready -> rsp_xbar_demux_022:src0_ready
	wire          rsp_xbar_demux_023_src0_endofpacket;                                                                // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_002:sink8_endofpacket
	wire          rsp_xbar_demux_023_src0_valid;                                                                      // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_002:sink8_valid
	wire          rsp_xbar_demux_023_src0_startofpacket;                                                              // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_002:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_023_src0_data;                                                                       // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_002:sink8_data
	wire   [54:0] rsp_xbar_demux_023_src0_channel;                                                                    // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_002:sink8_channel
	wire          rsp_xbar_demux_023_src0_ready;                                                                      // rsp_xbar_mux_002:sink8_ready -> rsp_xbar_demux_023:src0_ready
	wire          rsp_xbar_demux_023_src1_endofpacket;                                                                // rsp_xbar_demux_023:src1_endofpacket -> rsp_xbar_mux_003:sink2_endofpacket
	wire          rsp_xbar_demux_023_src1_valid;                                                                      // rsp_xbar_demux_023:src1_valid -> rsp_xbar_mux_003:sink2_valid
	wire          rsp_xbar_demux_023_src1_startofpacket;                                                              // rsp_xbar_demux_023:src1_startofpacket -> rsp_xbar_mux_003:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_023_src1_data;                                                                       // rsp_xbar_demux_023:src1_data -> rsp_xbar_mux_003:sink2_data
	wire   [54:0] rsp_xbar_demux_023_src1_channel;                                                                    // rsp_xbar_demux_023:src1_channel -> rsp_xbar_mux_003:sink2_channel
	wire          rsp_xbar_demux_023_src1_ready;                                                                      // rsp_xbar_mux_003:sink2_ready -> rsp_xbar_demux_023:src1_ready
	wire          rsp_xbar_demux_024_src0_endofpacket;                                                                // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_003:sink3_endofpacket
	wire          rsp_xbar_demux_024_src0_valid;                                                                      // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_003:sink3_valid
	wire          rsp_xbar_demux_024_src0_startofpacket;                                                              // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_003:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_024_src0_data;                                                                       // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_003:sink3_data
	wire   [54:0] rsp_xbar_demux_024_src0_channel;                                                                    // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_003:sink3_channel
	wire          rsp_xbar_demux_024_src0_ready;                                                                      // rsp_xbar_mux_003:sink3_ready -> rsp_xbar_demux_024:src0_ready
	wire          rsp_xbar_demux_024_src1_endofpacket;                                                                // rsp_xbar_demux_024:src1_endofpacket -> rsp_xbar_mux_008:sink2_endofpacket
	wire          rsp_xbar_demux_024_src1_valid;                                                                      // rsp_xbar_demux_024:src1_valid -> rsp_xbar_mux_008:sink2_valid
	wire          rsp_xbar_demux_024_src1_startofpacket;                                                              // rsp_xbar_demux_024:src1_startofpacket -> rsp_xbar_mux_008:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_024_src1_data;                                                                       // rsp_xbar_demux_024:src1_data -> rsp_xbar_mux_008:sink2_data
	wire   [54:0] rsp_xbar_demux_024_src1_channel;                                                                    // rsp_xbar_demux_024:src1_channel -> rsp_xbar_mux_008:sink2_channel
	wire          rsp_xbar_demux_024_src1_ready;                                                                      // rsp_xbar_mux_008:sink2_ready -> rsp_xbar_demux_024:src1_ready
	wire          rsp_xbar_demux_025_src0_endofpacket;                                                                // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_003:sink4_endofpacket
	wire          rsp_xbar_demux_025_src0_valid;                                                                      // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_003:sink4_valid
	wire          rsp_xbar_demux_025_src0_startofpacket;                                                              // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_003:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_025_src0_data;                                                                       // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_003:sink4_data
	wire   [54:0] rsp_xbar_demux_025_src0_channel;                                                                    // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_003:sink4_channel
	wire          rsp_xbar_demux_025_src0_ready;                                                                      // rsp_xbar_mux_003:sink4_ready -> rsp_xbar_demux_025:src0_ready
	wire          rsp_xbar_demux_025_src1_endofpacket;                                                                // rsp_xbar_demux_025:src1_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	wire          rsp_xbar_demux_025_src1_valid;                                                                      // rsp_xbar_demux_025:src1_valid -> rsp_xbar_mux_004:sink1_valid
	wire          rsp_xbar_demux_025_src1_startofpacket;                                                              // rsp_xbar_demux_025:src1_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_025_src1_data;                                                                       // rsp_xbar_demux_025:src1_data -> rsp_xbar_mux_004:sink1_data
	wire   [54:0] rsp_xbar_demux_025_src1_channel;                                                                    // rsp_xbar_demux_025:src1_channel -> rsp_xbar_mux_004:sink1_channel
	wire          rsp_xbar_demux_025_src1_ready;                                                                      // rsp_xbar_mux_004:sink1_ready -> rsp_xbar_demux_025:src1_ready
	wire          rsp_xbar_demux_026_src0_endofpacket;                                                                // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_003:sink5_endofpacket
	wire          rsp_xbar_demux_026_src0_valid;                                                                      // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_003:sink5_valid
	wire          rsp_xbar_demux_026_src0_startofpacket;                                                              // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_003:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_026_src0_data;                                                                       // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_003:sink5_data
	wire   [54:0] rsp_xbar_demux_026_src0_channel;                                                                    // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_003:sink5_channel
	wire          rsp_xbar_demux_026_src0_ready;                                                                      // rsp_xbar_mux_003:sink5_ready -> rsp_xbar_demux_026:src0_ready
	wire          rsp_xbar_demux_026_src1_endofpacket;                                                                // rsp_xbar_demux_026:src1_endofpacket -> rsp_xbar_mux_004:sink2_endofpacket
	wire          rsp_xbar_demux_026_src1_valid;                                                                      // rsp_xbar_demux_026:src1_valid -> rsp_xbar_mux_004:sink2_valid
	wire          rsp_xbar_demux_026_src1_startofpacket;                                                              // rsp_xbar_demux_026:src1_startofpacket -> rsp_xbar_mux_004:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_026_src1_data;                                                                       // rsp_xbar_demux_026:src1_data -> rsp_xbar_mux_004:sink2_data
	wire   [54:0] rsp_xbar_demux_026_src1_channel;                                                                    // rsp_xbar_demux_026:src1_channel -> rsp_xbar_mux_004:sink2_channel
	wire          rsp_xbar_demux_026_src1_ready;                                                                      // rsp_xbar_mux_004:sink2_ready -> rsp_xbar_demux_026:src1_ready
	wire          rsp_xbar_demux_027_src0_endofpacket;                                                                // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_003:sink6_endofpacket
	wire          rsp_xbar_demux_027_src0_valid;                                                                      // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_003:sink6_valid
	wire          rsp_xbar_demux_027_src0_startofpacket;                                                              // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_003:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_027_src0_data;                                                                       // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_003:sink6_data
	wire   [54:0] rsp_xbar_demux_027_src0_channel;                                                                    // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_003:sink6_channel
	wire          rsp_xbar_demux_027_src0_ready;                                                                      // rsp_xbar_mux_003:sink6_ready -> rsp_xbar_demux_027:src0_ready
	wire          rsp_xbar_demux_028_src0_endofpacket;                                                                // rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux_003:sink7_endofpacket
	wire          rsp_xbar_demux_028_src0_valid;                                                                      // rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux_003:sink7_valid
	wire          rsp_xbar_demux_028_src0_startofpacket;                                                              // rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux_003:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_028_src0_data;                                                                       // rsp_xbar_demux_028:src0_data -> rsp_xbar_mux_003:sink7_data
	wire   [54:0] rsp_xbar_demux_028_src0_channel;                                                                    // rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux_003:sink7_channel
	wire          rsp_xbar_demux_028_src0_ready;                                                                      // rsp_xbar_mux_003:sink7_ready -> rsp_xbar_demux_028:src0_ready
	wire          rsp_xbar_demux_029_src0_endofpacket;                                                                // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_003:sink8_endofpacket
	wire          rsp_xbar_demux_029_src0_valid;                                                                      // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_003:sink8_valid
	wire          rsp_xbar_demux_029_src0_startofpacket;                                                              // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_003:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_029_src0_data;                                                                       // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_003:sink8_data
	wire   [54:0] rsp_xbar_demux_029_src0_channel;                                                                    // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_003:sink8_channel
	wire          rsp_xbar_demux_029_src0_ready;                                                                      // rsp_xbar_mux_003:sink8_ready -> rsp_xbar_demux_029:src0_ready
	wire          rsp_xbar_demux_030_src0_endofpacket;                                                                // rsp_xbar_demux_030:src0_endofpacket -> rsp_xbar_mux_003:sink9_endofpacket
	wire          rsp_xbar_demux_030_src0_valid;                                                                      // rsp_xbar_demux_030:src0_valid -> rsp_xbar_mux_003:sink9_valid
	wire          rsp_xbar_demux_030_src0_startofpacket;                                                              // rsp_xbar_demux_030:src0_startofpacket -> rsp_xbar_mux_003:sink9_startofpacket
	wire  [106:0] rsp_xbar_demux_030_src0_data;                                                                       // rsp_xbar_demux_030:src0_data -> rsp_xbar_mux_003:sink9_data
	wire   [54:0] rsp_xbar_demux_030_src0_channel;                                                                    // rsp_xbar_demux_030:src0_channel -> rsp_xbar_mux_003:sink9_channel
	wire          rsp_xbar_demux_030_src0_ready;                                                                      // rsp_xbar_mux_003:sink9_ready -> rsp_xbar_demux_030:src0_ready
	wire          rsp_xbar_demux_031_src0_endofpacket;                                                                // rsp_xbar_demux_031:src0_endofpacket -> rsp_xbar_mux_003:sink10_endofpacket
	wire          rsp_xbar_demux_031_src0_valid;                                                                      // rsp_xbar_demux_031:src0_valid -> rsp_xbar_mux_003:sink10_valid
	wire          rsp_xbar_demux_031_src0_startofpacket;                                                              // rsp_xbar_demux_031:src0_startofpacket -> rsp_xbar_mux_003:sink10_startofpacket
	wire  [106:0] rsp_xbar_demux_031_src0_data;                                                                       // rsp_xbar_demux_031:src0_data -> rsp_xbar_mux_003:sink10_data
	wire   [54:0] rsp_xbar_demux_031_src0_channel;                                                                    // rsp_xbar_demux_031:src0_channel -> rsp_xbar_mux_003:sink10_channel
	wire          rsp_xbar_demux_031_src0_ready;                                                                      // rsp_xbar_mux_003:sink10_ready -> rsp_xbar_demux_031:src0_ready
	wire          rsp_xbar_demux_032_src0_endofpacket;                                                                // rsp_xbar_demux_032:src0_endofpacket -> rsp_xbar_mux_005:sink1_endofpacket
	wire          rsp_xbar_demux_032_src0_valid;                                                                      // rsp_xbar_demux_032:src0_valid -> rsp_xbar_mux_005:sink1_valid
	wire          rsp_xbar_demux_032_src0_startofpacket;                                                              // rsp_xbar_demux_032:src0_startofpacket -> rsp_xbar_mux_005:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_032_src0_data;                                                                       // rsp_xbar_demux_032:src0_data -> rsp_xbar_mux_005:sink1_data
	wire   [54:0] rsp_xbar_demux_032_src0_channel;                                                                    // rsp_xbar_demux_032:src0_channel -> rsp_xbar_mux_005:sink1_channel
	wire          rsp_xbar_demux_032_src0_ready;                                                                      // rsp_xbar_mux_005:sink1_ready -> rsp_xbar_demux_032:src0_ready
	wire          rsp_xbar_demux_032_src1_endofpacket;                                                                // rsp_xbar_demux_032:src1_endofpacket -> rsp_xbar_mux_006:sink4_endofpacket
	wire          rsp_xbar_demux_032_src1_valid;                                                                      // rsp_xbar_demux_032:src1_valid -> rsp_xbar_mux_006:sink4_valid
	wire          rsp_xbar_demux_032_src1_startofpacket;                                                              // rsp_xbar_demux_032:src1_startofpacket -> rsp_xbar_mux_006:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_032_src1_data;                                                                       // rsp_xbar_demux_032:src1_data -> rsp_xbar_mux_006:sink4_data
	wire   [54:0] rsp_xbar_demux_032_src1_channel;                                                                    // rsp_xbar_demux_032:src1_channel -> rsp_xbar_mux_006:sink4_channel
	wire          rsp_xbar_demux_032_src1_ready;                                                                      // rsp_xbar_mux_006:sink4_ready -> rsp_xbar_demux_032:src1_ready
	wire          rsp_xbar_demux_033_src0_endofpacket;                                                                // rsp_xbar_demux_033:src0_endofpacket -> rsp_xbar_mux_005:sink2_endofpacket
	wire          rsp_xbar_demux_033_src0_valid;                                                                      // rsp_xbar_demux_033:src0_valid -> rsp_xbar_mux_005:sink2_valid
	wire          rsp_xbar_demux_033_src0_startofpacket;                                                              // rsp_xbar_demux_033:src0_startofpacket -> rsp_xbar_mux_005:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_033_src0_data;                                                                       // rsp_xbar_demux_033:src0_data -> rsp_xbar_mux_005:sink2_data
	wire   [54:0] rsp_xbar_demux_033_src0_channel;                                                                    // rsp_xbar_demux_033:src0_channel -> rsp_xbar_mux_005:sink2_channel
	wire          rsp_xbar_demux_033_src0_ready;                                                                      // rsp_xbar_mux_005:sink2_ready -> rsp_xbar_demux_033:src0_ready
	wire          rsp_xbar_demux_033_src1_endofpacket;                                                                // rsp_xbar_demux_033:src1_endofpacket -> rsp_xbar_mux_006:sink5_endofpacket
	wire          rsp_xbar_demux_033_src1_valid;                                                                      // rsp_xbar_demux_033:src1_valid -> rsp_xbar_mux_006:sink5_valid
	wire          rsp_xbar_demux_033_src1_startofpacket;                                                              // rsp_xbar_demux_033:src1_startofpacket -> rsp_xbar_mux_006:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_033_src1_data;                                                                       // rsp_xbar_demux_033:src1_data -> rsp_xbar_mux_006:sink5_data
	wire   [54:0] rsp_xbar_demux_033_src1_channel;                                                                    // rsp_xbar_demux_033:src1_channel -> rsp_xbar_mux_006:sink5_channel
	wire          rsp_xbar_demux_033_src1_ready;                                                                      // rsp_xbar_mux_006:sink5_ready -> rsp_xbar_demux_033:src1_ready
	wire          rsp_xbar_demux_034_src0_endofpacket;                                                                // rsp_xbar_demux_034:src0_endofpacket -> rsp_xbar_mux_006:sink6_endofpacket
	wire          rsp_xbar_demux_034_src0_valid;                                                                      // rsp_xbar_demux_034:src0_valid -> rsp_xbar_mux_006:sink6_valid
	wire          rsp_xbar_demux_034_src0_startofpacket;                                                              // rsp_xbar_demux_034:src0_startofpacket -> rsp_xbar_mux_006:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_034_src0_data;                                                                       // rsp_xbar_demux_034:src0_data -> rsp_xbar_mux_006:sink6_data
	wire   [54:0] rsp_xbar_demux_034_src0_channel;                                                                    // rsp_xbar_demux_034:src0_channel -> rsp_xbar_mux_006:sink6_channel
	wire          rsp_xbar_demux_034_src0_ready;                                                                      // rsp_xbar_mux_006:sink6_ready -> rsp_xbar_demux_034:src0_ready
	wire          rsp_xbar_demux_035_src0_endofpacket;                                                                // rsp_xbar_demux_035:src0_endofpacket -> rsp_xbar_mux_006:sink7_endofpacket
	wire          rsp_xbar_demux_035_src0_valid;                                                                      // rsp_xbar_demux_035:src0_valid -> rsp_xbar_mux_006:sink7_valid
	wire          rsp_xbar_demux_035_src0_startofpacket;                                                              // rsp_xbar_demux_035:src0_startofpacket -> rsp_xbar_mux_006:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_035_src0_data;                                                                       // rsp_xbar_demux_035:src0_data -> rsp_xbar_mux_006:sink7_data
	wire   [54:0] rsp_xbar_demux_035_src0_channel;                                                                    // rsp_xbar_demux_035:src0_channel -> rsp_xbar_mux_006:sink7_channel
	wire          rsp_xbar_demux_035_src0_ready;                                                                      // rsp_xbar_mux_006:sink7_ready -> rsp_xbar_demux_035:src0_ready
	wire          rsp_xbar_demux_036_src0_endofpacket;                                                                // rsp_xbar_demux_036:src0_endofpacket -> rsp_xbar_mux_006:sink8_endofpacket
	wire          rsp_xbar_demux_036_src0_valid;                                                                      // rsp_xbar_demux_036:src0_valid -> rsp_xbar_mux_006:sink8_valid
	wire          rsp_xbar_demux_036_src0_startofpacket;                                                              // rsp_xbar_demux_036:src0_startofpacket -> rsp_xbar_mux_006:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_036_src0_data;                                                                       // rsp_xbar_demux_036:src0_data -> rsp_xbar_mux_006:sink8_data
	wire   [54:0] rsp_xbar_demux_036_src0_channel;                                                                    // rsp_xbar_demux_036:src0_channel -> rsp_xbar_mux_006:sink8_channel
	wire          rsp_xbar_demux_036_src0_ready;                                                                      // rsp_xbar_mux_006:sink8_ready -> rsp_xbar_demux_036:src0_ready
	wire          rsp_xbar_demux_037_src0_endofpacket;                                                                // rsp_xbar_demux_037:src0_endofpacket -> rsp_xbar_mux_006:sink9_endofpacket
	wire          rsp_xbar_demux_037_src0_valid;                                                                      // rsp_xbar_demux_037:src0_valid -> rsp_xbar_mux_006:sink9_valid
	wire          rsp_xbar_demux_037_src0_startofpacket;                                                              // rsp_xbar_demux_037:src0_startofpacket -> rsp_xbar_mux_006:sink9_startofpacket
	wire  [106:0] rsp_xbar_demux_037_src0_data;                                                                       // rsp_xbar_demux_037:src0_data -> rsp_xbar_mux_006:sink9_data
	wire   [54:0] rsp_xbar_demux_037_src0_channel;                                                                    // rsp_xbar_demux_037:src0_channel -> rsp_xbar_mux_006:sink9_channel
	wire          rsp_xbar_demux_037_src0_ready;                                                                      // rsp_xbar_mux_006:sink9_ready -> rsp_xbar_demux_037:src0_ready
	wire          rsp_xbar_demux_038_src0_endofpacket;                                                                // rsp_xbar_demux_038:src0_endofpacket -> rsp_xbar_mux_006:sink10_endofpacket
	wire          rsp_xbar_demux_038_src0_valid;                                                                      // rsp_xbar_demux_038:src0_valid -> rsp_xbar_mux_006:sink10_valid
	wire          rsp_xbar_demux_038_src0_startofpacket;                                                              // rsp_xbar_demux_038:src0_startofpacket -> rsp_xbar_mux_006:sink10_startofpacket
	wire  [106:0] rsp_xbar_demux_038_src0_data;                                                                       // rsp_xbar_demux_038:src0_data -> rsp_xbar_mux_006:sink10_data
	wire   [54:0] rsp_xbar_demux_038_src0_channel;                                                                    // rsp_xbar_demux_038:src0_channel -> rsp_xbar_mux_006:sink10_channel
	wire          rsp_xbar_demux_038_src0_ready;                                                                      // rsp_xbar_mux_006:sink10_ready -> rsp_xbar_demux_038:src0_ready
	wire          rsp_xbar_demux_039_src0_endofpacket;                                                                // rsp_xbar_demux_039:src0_endofpacket -> rsp_xbar_mux_006:sink11_endofpacket
	wire          rsp_xbar_demux_039_src0_valid;                                                                      // rsp_xbar_demux_039:src0_valid -> rsp_xbar_mux_006:sink11_valid
	wire          rsp_xbar_demux_039_src0_startofpacket;                                                              // rsp_xbar_demux_039:src0_startofpacket -> rsp_xbar_mux_006:sink11_startofpacket
	wire  [106:0] rsp_xbar_demux_039_src0_data;                                                                       // rsp_xbar_demux_039:src0_data -> rsp_xbar_mux_006:sink11_data
	wire   [54:0] rsp_xbar_demux_039_src0_channel;                                                                    // rsp_xbar_demux_039:src0_channel -> rsp_xbar_mux_006:sink11_channel
	wire          rsp_xbar_demux_039_src0_ready;                                                                      // rsp_xbar_mux_006:sink11_ready -> rsp_xbar_demux_039:src0_ready
	wire          rsp_xbar_demux_040_src0_endofpacket;                                                                // rsp_xbar_demux_040:src0_endofpacket -> rsp_xbar_mux_006:sink12_endofpacket
	wire          rsp_xbar_demux_040_src0_valid;                                                                      // rsp_xbar_demux_040:src0_valid -> rsp_xbar_mux_006:sink12_valid
	wire          rsp_xbar_demux_040_src0_startofpacket;                                                              // rsp_xbar_demux_040:src0_startofpacket -> rsp_xbar_mux_006:sink12_startofpacket
	wire  [106:0] rsp_xbar_demux_040_src0_data;                                                                       // rsp_xbar_demux_040:src0_data -> rsp_xbar_mux_006:sink12_data
	wire   [54:0] rsp_xbar_demux_040_src0_channel;                                                                    // rsp_xbar_demux_040:src0_channel -> rsp_xbar_mux_006:sink12_channel
	wire          rsp_xbar_demux_040_src0_ready;                                                                      // rsp_xbar_mux_006:sink12_ready -> rsp_xbar_demux_040:src0_ready
	wire          rsp_xbar_demux_040_src1_endofpacket;                                                                // rsp_xbar_demux_040:src1_endofpacket -> rsp_xbar_mux_007:sink1_endofpacket
	wire          rsp_xbar_demux_040_src1_valid;                                                                      // rsp_xbar_demux_040:src1_valid -> rsp_xbar_mux_007:sink1_valid
	wire          rsp_xbar_demux_040_src1_startofpacket;                                                              // rsp_xbar_demux_040:src1_startofpacket -> rsp_xbar_mux_007:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_040_src1_data;                                                                       // rsp_xbar_demux_040:src1_data -> rsp_xbar_mux_007:sink1_data
	wire   [54:0] rsp_xbar_demux_040_src1_channel;                                                                    // rsp_xbar_demux_040:src1_channel -> rsp_xbar_mux_007:sink1_channel
	wire          rsp_xbar_demux_040_src1_ready;                                                                      // rsp_xbar_mux_007:sink1_ready -> rsp_xbar_demux_040:src1_ready
	wire          rsp_xbar_demux_041_src0_endofpacket;                                                                // rsp_xbar_demux_041:src0_endofpacket -> rsp_xbar_mux_007:sink2_endofpacket
	wire          rsp_xbar_demux_041_src0_valid;                                                                      // rsp_xbar_demux_041:src0_valid -> rsp_xbar_mux_007:sink2_valid
	wire          rsp_xbar_demux_041_src0_startofpacket;                                                              // rsp_xbar_demux_041:src0_startofpacket -> rsp_xbar_mux_007:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_041_src0_data;                                                                       // rsp_xbar_demux_041:src0_data -> rsp_xbar_mux_007:sink2_data
	wire   [54:0] rsp_xbar_demux_041_src0_channel;                                                                    // rsp_xbar_demux_041:src0_channel -> rsp_xbar_mux_007:sink2_channel
	wire          rsp_xbar_demux_041_src0_ready;                                                                      // rsp_xbar_mux_007:sink2_ready -> rsp_xbar_demux_041:src0_ready
	wire          rsp_xbar_demux_041_src1_endofpacket;                                                                // rsp_xbar_demux_041:src1_endofpacket -> rsp_xbar_mux_010:sink1_endofpacket
	wire          rsp_xbar_demux_041_src1_valid;                                                                      // rsp_xbar_demux_041:src1_valid -> rsp_xbar_mux_010:sink1_valid
	wire          rsp_xbar_demux_041_src1_startofpacket;                                                              // rsp_xbar_demux_041:src1_startofpacket -> rsp_xbar_mux_010:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_041_src1_data;                                                                       // rsp_xbar_demux_041:src1_data -> rsp_xbar_mux_010:sink1_data
	wire   [54:0] rsp_xbar_demux_041_src1_channel;                                                                    // rsp_xbar_demux_041:src1_channel -> rsp_xbar_mux_010:sink1_channel
	wire          rsp_xbar_demux_041_src1_ready;                                                                      // rsp_xbar_mux_010:sink1_ready -> rsp_xbar_demux_041:src1_ready
	wire          rsp_xbar_demux_042_src0_endofpacket;                                                                // rsp_xbar_demux_042:src0_endofpacket -> rsp_xbar_mux_007:sink3_endofpacket
	wire          rsp_xbar_demux_042_src0_valid;                                                                      // rsp_xbar_demux_042:src0_valid -> rsp_xbar_mux_007:sink3_valid
	wire          rsp_xbar_demux_042_src0_startofpacket;                                                              // rsp_xbar_demux_042:src0_startofpacket -> rsp_xbar_mux_007:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_042_src0_data;                                                                       // rsp_xbar_demux_042:src0_data -> rsp_xbar_mux_007:sink3_data
	wire   [54:0] rsp_xbar_demux_042_src0_channel;                                                                    // rsp_xbar_demux_042:src0_channel -> rsp_xbar_mux_007:sink3_channel
	wire          rsp_xbar_demux_042_src0_ready;                                                                      // rsp_xbar_mux_007:sink3_ready -> rsp_xbar_demux_042:src0_ready
	wire          rsp_xbar_demux_042_src1_endofpacket;                                                                // rsp_xbar_demux_042:src1_endofpacket -> rsp_xbar_mux_010:sink2_endofpacket
	wire          rsp_xbar_demux_042_src1_valid;                                                                      // rsp_xbar_demux_042:src1_valid -> rsp_xbar_mux_010:sink2_valid
	wire          rsp_xbar_demux_042_src1_startofpacket;                                                              // rsp_xbar_demux_042:src1_startofpacket -> rsp_xbar_mux_010:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_042_src1_data;                                                                       // rsp_xbar_demux_042:src1_data -> rsp_xbar_mux_010:sink2_data
	wire   [54:0] rsp_xbar_demux_042_src1_channel;                                                                    // rsp_xbar_demux_042:src1_channel -> rsp_xbar_mux_010:sink2_channel
	wire          rsp_xbar_demux_042_src1_ready;                                                                      // rsp_xbar_mux_010:sink2_ready -> rsp_xbar_demux_042:src1_ready
	wire          rsp_xbar_demux_043_src0_endofpacket;                                                                // rsp_xbar_demux_043:src0_endofpacket -> rsp_xbar_mux_007:sink4_endofpacket
	wire          rsp_xbar_demux_043_src0_valid;                                                                      // rsp_xbar_demux_043:src0_valid -> rsp_xbar_mux_007:sink4_valid
	wire          rsp_xbar_demux_043_src0_startofpacket;                                                              // rsp_xbar_demux_043:src0_startofpacket -> rsp_xbar_mux_007:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_043_src0_data;                                                                       // rsp_xbar_demux_043:src0_data -> rsp_xbar_mux_007:sink4_data
	wire   [54:0] rsp_xbar_demux_043_src0_channel;                                                                    // rsp_xbar_demux_043:src0_channel -> rsp_xbar_mux_007:sink4_channel
	wire          rsp_xbar_demux_043_src0_ready;                                                                      // rsp_xbar_mux_007:sink4_ready -> rsp_xbar_demux_043:src0_ready
	wire          rsp_xbar_demux_044_src0_endofpacket;                                                                // rsp_xbar_demux_044:src0_endofpacket -> rsp_xbar_mux_007:sink5_endofpacket
	wire          rsp_xbar_demux_044_src0_valid;                                                                      // rsp_xbar_demux_044:src0_valid -> rsp_xbar_mux_007:sink5_valid
	wire          rsp_xbar_demux_044_src0_startofpacket;                                                              // rsp_xbar_demux_044:src0_startofpacket -> rsp_xbar_mux_007:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_044_src0_data;                                                                       // rsp_xbar_demux_044:src0_data -> rsp_xbar_mux_007:sink5_data
	wire   [54:0] rsp_xbar_demux_044_src0_channel;                                                                    // rsp_xbar_demux_044:src0_channel -> rsp_xbar_mux_007:sink5_channel
	wire          rsp_xbar_demux_044_src0_ready;                                                                      // rsp_xbar_mux_007:sink5_ready -> rsp_xbar_demux_044:src0_ready
	wire          rsp_xbar_demux_045_src0_endofpacket;                                                                // rsp_xbar_demux_045:src0_endofpacket -> rsp_xbar_mux_007:sink6_endofpacket
	wire          rsp_xbar_demux_045_src0_valid;                                                                      // rsp_xbar_demux_045:src0_valid -> rsp_xbar_mux_007:sink6_valid
	wire          rsp_xbar_demux_045_src0_startofpacket;                                                              // rsp_xbar_demux_045:src0_startofpacket -> rsp_xbar_mux_007:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_045_src0_data;                                                                       // rsp_xbar_demux_045:src0_data -> rsp_xbar_mux_007:sink6_data
	wire   [54:0] rsp_xbar_demux_045_src0_channel;                                                                    // rsp_xbar_demux_045:src0_channel -> rsp_xbar_mux_007:sink6_channel
	wire          rsp_xbar_demux_045_src0_ready;                                                                      // rsp_xbar_mux_007:sink6_ready -> rsp_xbar_demux_045:src0_ready
	wire          rsp_xbar_demux_046_src0_endofpacket;                                                                // rsp_xbar_demux_046:src0_endofpacket -> rsp_xbar_mux_007:sink7_endofpacket
	wire          rsp_xbar_demux_046_src0_valid;                                                                      // rsp_xbar_demux_046:src0_valid -> rsp_xbar_mux_007:sink7_valid
	wire          rsp_xbar_demux_046_src0_startofpacket;                                                              // rsp_xbar_demux_046:src0_startofpacket -> rsp_xbar_mux_007:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_046_src0_data;                                                                       // rsp_xbar_demux_046:src0_data -> rsp_xbar_mux_007:sink7_data
	wire   [54:0] rsp_xbar_demux_046_src0_channel;                                                                    // rsp_xbar_demux_046:src0_channel -> rsp_xbar_mux_007:sink7_channel
	wire          rsp_xbar_demux_046_src0_ready;                                                                      // rsp_xbar_mux_007:sink7_ready -> rsp_xbar_demux_046:src0_ready
	wire          rsp_xbar_demux_047_src0_endofpacket;                                                                // rsp_xbar_demux_047:src0_endofpacket -> rsp_xbar_mux_007:sink8_endofpacket
	wire          rsp_xbar_demux_047_src0_valid;                                                                      // rsp_xbar_demux_047:src0_valid -> rsp_xbar_mux_007:sink8_valid
	wire          rsp_xbar_demux_047_src0_startofpacket;                                                              // rsp_xbar_demux_047:src0_startofpacket -> rsp_xbar_mux_007:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_047_src0_data;                                                                       // rsp_xbar_demux_047:src0_data -> rsp_xbar_mux_007:sink8_data
	wire   [54:0] rsp_xbar_demux_047_src0_channel;                                                                    // rsp_xbar_demux_047:src0_channel -> rsp_xbar_mux_007:sink8_channel
	wire          rsp_xbar_demux_047_src0_ready;                                                                      // rsp_xbar_mux_007:sink8_ready -> rsp_xbar_demux_047:src0_ready
	wire          rsp_xbar_demux_047_src1_endofpacket;                                                                // rsp_xbar_demux_047:src1_endofpacket -> rsp_xbar_mux_008:sink3_endofpacket
	wire          rsp_xbar_demux_047_src1_valid;                                                                      // rsp_xbar_demux_047:src1_valid -> rsp_xbar_mux_008:sink3_valid
	wire          rsp_xbar_demux_047_src1_startofpacket;                                                              // rsp_xbar_demux_047:src1_startofpacket -> rsp_xbar_mux_008:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_047_src1_data;                                                                       // rsp_xbar_demux_047:src1_data -> rsp_xbar_mux_008:sink3_data
	wire   [54:0] rsp_xbar_demux_047_src1_channel;                                                                    // rsp_xbar_demux_047:src1_channel -> rsp_xbar_mux_008:sink3_channel
	wire          rsp_xbar_demux_047_src1_ready;                                                                      // rsp_xbar_mux_008:sink3_ready -> rsp_xbar_demux_047:src1_ready
	wire          rsp_xbar_demux_048_src0_endofpacket;                                                                // rsp_xbar_demux_048:src0_endofpacket -> rsp_xbar_mux_008:sink4_endofpacket
	wire          rsp_xbar_demux_048_src0_valid;                                                                      // rsp_xbar_demux_048:src0_valid -> rsp_xbar_mux_008:sink4_valid
	wire          rsp_xbar_demux_048_src0_startofpacket;                                                              // rsp_xbar_demux_048:src0_startofpacket -> rsp_xbar_mux_008:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_048_src0_data;                                                                       // rsp_xbar_demux_048:src0_data -> rsp_xbar_mux_008:sink4_data
	wire   [54:0] rsp_xbar_demux_048_src0_channel;                                                                    // rsp_xbar_demux_048:src0_channel -> rsp_xbar_mux_008:sink4_channel
	wire          rsp_xbar_demux_048_src0_ready;                                                                      // rsp_xbar_mux_008:sink4_ready -> rsp_xbar_demux_048:src0_ready
	wire          rsp_xbar_demux_048_src1_endofpacket;                                                                // rsp_xbar_demux_048:src1_endofpacket -> rsp_xbar_mux_009:sink1_endofpacket
	wire          rsp_xbar_demux_048_src1_valid;                                                                      // rsp_xbar_demux_048:src1_valid -> rsp_xbar_mux_009:sink1_valid
	wire          rsp_xbar_demux_048_src1_startofpacket;                                                              // rsp_xbar_demux_048:src1_startofpacket -> rsp_xbar_mux_009:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_048_src1_data;                                                                       // rsp_xbar_demux_048:src1_data -> rsp_xbar_mux_009:sink1_data
	wire   [54:0] rsp_xbar_demux_048_src1_channel;                                                                    // rsp_xbar_demux_048:src1_channel -> rsp_xbar_mux_009:sink1_channel
	wire          rsp_xbar_demux_048_src1_ready;                                                                      // rsp_xbar_mux_009:sink1_ready -> rsp_xbar_demux_048:src1_ready
	wire          rsp_xbar_demux_049_src0_endofpacket;                                                                // rsp_xbar_demux_049:src0_endofpacket -> rsp_xbar_mux_008:sink5_endofpacket
	wire          rsp_xbar_demux_049_src0_valid;                                                                      // rsp_xbar_demux_049:src0_valid -> rsp_xbar_mux_008:sink5_valid
	wire          rsp_xbar_demux_049_src0_startofpacket;                                                              // rsp_xbar_demux_049:src0_startofpacket -> rsp_xbar_mux_008:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_049_src0_data;                                                                       // rsp_xbar_demux_049:src0_data -> rsp_xbar_mux_008:sink5_data
	wire   [54:0] rsp_xbar_demux_049_src0_channel;                                                                    // rsp_xbar_demux_049:src0_channel -> rsp_xbar_mux_008:sink5_channel
	wire          rsp_xbar_demux_049_src0_ready;                                                                      // rsp_xbar_mux_008:sink5_ready -> rsp_xbar_demux_049:src0_ready
	wire          rsp_xbar_demux_049_src1_endofpacket;                                                                // rsp_xbar_demux_049:src1_endofpacket -> rsp_xbar_mux_009:sink2_endofpacket
	wire          rsp_xbar_demux_049_src1_valid;                                                                      // rsp_xbar_demux_049:src1_valid -> rsp_xbar_mux_009:sink2_valid
	wire          rsp_xbar_demux_049_src1_startofpacket;                                                              // rsp_xbar_demux_049:src1_startofpacket -> rsp_xbar_mux_009:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_049_src1_data;                                                                       // rsp_xbar_demux_049:src1_data -> rsp_xbar_mux_009:sink2_data
	wire   [54:0] rsp_xbar_demux_049_src1_channel;                                                                    // rsp_xbar_demux_049:src1_channel -> rsp_xbar_mux_009:sink2_channel
	wire          rsp_xbar_demux_049_src1_ready;                                                                      // rsp_xbar_mux_009:sink2_ready -> rsp_xbar_demux_049:src1_ready
	wire          rsp_xbar_demux_050_src0_endofpacket;                                                                // rsp_xbar_demux_050:src0_endofpacket -> rsp_xbar_mux_008:sink6_endofpacket
	wire          rsp_xbar_demux_050_src0_valid;                                                                      // rsp_xbar_demux_050:src0_valid -> rsp_xbar_mux_008:sink6_valid
	wire          rsp_xbar_demux_050_src0_startofpacket;                                                              // rsp_xbar_demux_050:src0_startofpacket -> rsp_xbar_mux_008:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_050_src0_data;                                                                       // rsp_xbar_demux_050:src0_data -> rsp_xbar_mux_008:sink6_data
	wire   [54:0] rsp_xbar_demux_050_src0_channel;                                                                    // rsp_xbar_demux_050:src0_channel -> rsp_xbar_mux_008:sink6_channel
	wire          rsp_xbar_demux_050_src0_ready;                                                                      // rsp_xbar_mux_008:sink6_ready -> rsp_xbar_demux_050:src0_ready
	wire          rsp_xbar_demux_051_src0_endofpacket;                                                                // rsp_xbar_demux_051:src0_endofpacket -> rsp_xbar_mux_008:sink7_endofpacket
	wire          rsp_xbar_demux_051_src0_valid;                                                                      // rsp_xbar_demux_051:src0_valid -> rsp_xbar_mux_008:sink7_valid
	wire          rsp_xbar_demux_051_src0_startofpacket;                                                              // rsp_xbar_demux_051:src0_startofpacket -> rsp_xbar_mux_008:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_051_src0_data;                                                                       // rsp_xbar_demux_051:src0_data -> rsp_xbar_mux_008:sink7_data
	wire   [54:0] rsp_xbar_demux_051_src0_channel;                                                                    // rsp_xbar_demux_051:src0_channel -> rsp_xbar_mux_008:sink7_channel
	wire          rsp_xbar_demux_051_src0_ready;                                                                      // rsp_xbar_mux_008:sink7_ready -> rsp_xbar_demux_051:src0_ready
	wire          rsp_xbar_demux_052_src0_endofpacket;                                                                // rsp_xbar_demux_052:src0_endofpacket -> rsp_xbar_mux_008:sink8_endofpacket
	wire          rsp_xbar_demux_052_src0_valid;                                                                      // rsp_xbar_demux_052:src0_valid -> rsp_xbar_mux_008:sink8_valid
	wire          rsp_xbar_demux_052_src0_startofpacket;                                                              // rsp_xbar_demux_052:src0_startofpacket -> rsp_xbar_mux_008:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_052_src0_data;                                                                       // rsp_xbar_demux_052:src0_data -> rsp_xbar_mux_008:sink8_data
	wire   [54:0] rsp_xbar_demux_052_src0_channel;                                                                    // rsp_xbar_demux_052:src0_channel -> rsp_xbar_mux_008:sink8_channel
	wire          rsp_xbar_demux_052_src0_ready;                                                                      // rsp_xbar_mux_008:sink8_ready -> rsp_xbar_demux_052:src0_ready
	wire          rsp_xbar_demux_053_src0_endofpacket;                                                                // rsp_xbar_demux_053:src0_endofpacket -> rsp_xbar_mux_008:sink9_endofpacket
	wire          rsp_xbar_demux_053_src0_valid;                                                                      // rsp_xbar_demux_053:src0_valid -> rsp_xbar_mux_008:sink9_valid
	wire          rsp_xbar_demux_053_src0_startofpacket;                                                              // rsp_xbar_demux_053:src0_startofpacket -> rsp_xbar_mux_008:sink9_startofpacket
	wire  [106:0] rsp_xbar_demux_053_src0_data;                                                                       // rsp_xbar_demux_053:src0_data -> rsp_xbar_mux_008:sink9_data
	wire   [54:0] rsp_xbar_demux_053_src0_channel;                                                                    // rsp_xbar_demux_053:src0_channel -> rsp_xbar_mux_008:sink9_channel
	wire          rsp_xbar_demux_053_src0_ready;                                                                      // rsp_xbar_mux_008:sink9_ready -> rsp_xbar_demux_053:src0_ready
	wire          rsp_xbar_demux_054_src0_endofpacket;                                                                // rsp_xbar_demux_054:src0_endofpacket -> rsp_xbar_mux_008:sink10_endofpacket
	wire          rsp_xbar_demux_054_src0_valid;                                                                      // rsp_xbar_demux_054:src0_valid -> rsp_xbar_mux_008:sink10_valid
	wire          rsp_xbar_demux_054_src0_startofpacket;                                                              // rsp_xbar_demux_054:src0_startofpacket -> rsp_xbar_mux_008:sink10_startofpacket
	wire  [106:0] rsp_xbar_demux_054_src0_data;                                                                       // rsp_xbar_demux_054:src0_data -> rsp_xbar_mux_008:sink10_data
	wire   [54:0] rsp_xbar_demux_054_src0_channel;                                                                    // rsp_xbar_demux_054:src0_channel -> rsp_xbar_mux_008:sink10_channel
	wire          rsp_xbar_demux_054_src0_ready;                                                                      // rsp_xbar_mux_008:sink10_ready -> rsp_xbar_demux_054:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                        // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                      // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [106:0] limiter_cmd_src_data;                                                                               // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [54:0] limiter_cmd_src_channel;                                                                            // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                              // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                       // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                             // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                     // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_src_data;                                                                              // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [54:0] rsp_xbar_mux_src_channel;                                                                           // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                             // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                    // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                          // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                  // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [106:0] addr_router_001_src_data;                                                                           // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [54:0] addr_router_001_src_channel;                                                                        // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                          // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                   // rsp_xbar_mux_001:src_endofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                         // rsp_xbar_mux_001:src_valid -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                 // rsp_xbar_mux_001:src_startofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_001_src_data;                                                                          // rsp_xbar_mux_001:src_data -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] rsp_xbar_mux_001_src_channel;                                                                       // rsp_xbar_mux_001:src_channel -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                         // cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                    // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                          // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                  // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [106:0] addr_router_002_src_data;                                                                           // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [54:0] addr_router_002_src_channel;                                                                        // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                          // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                   // rsp_xbar_mux_002:src_endofpacket -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                         // rsp_xbar_mux_002:src_valid -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                                 // rsp_xbar_mux_002:src_startofpacket -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_002_src_data;                                                                          // rsp_xbar_mux_002:src_data -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] rsp_xbar_mux_002_src_channel;                                                                       // rsp_xbar_mux_002:src_channel -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                         // cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	wire          addr_router_003_src_endofpacket;                                                                    // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                          // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                  // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [106:0] addr_router_003_src_data;                                                                           // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire   [54:0] addr_router_003_src_channel;                                                                        // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                          // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                   // rsp_xbar_mux_003:src_endofpacket -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                         // rsp_xbar_mux_003:src_valid -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                                 // rsp_xbar_mux_003:src_startofpacket -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_003_src_data;                                                                          // rsp_xbar_mux_003:src_data -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] rsp_xbar_mux_003_src_channel;                                                                       // rsp_xbar_mux_003:src_channel -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                         // cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_003:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                    // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                  // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [106:0] limiter_001_cmd_src_data;                                                                           // limiter_001:cmd_src_data -> cmd_xbar_demux_004:sink_data
	wire   [54:0] limiter_001_cmd_src_channel;                                                                        // limiter_001:cmd_src_channel -> cmd_xbar_demux_004:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                          // cmd_xbar_demux_004:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_004_src_endofpacket;                                                                   // rsp_xbar_mux_004:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_004_src_valid;                                                                         // rsp_xbar_mux_004:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_004_src_startofpacket;                                                                 // rsp_xbar_mux_004:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_004_src_data;                                                                          // rsp_xbar_mux_004:src_data -> limiter_001:rsp_sink_data
	wire   [54:0] rsp_xbar_mux_004_src_channel;                                                                       // rsp_xbar_mux_004:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_004_src_ready;                                                                         // limiter_001:rsp_sink_ready -> rsp_xbar_mux_004:src_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                    // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                  // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [106:0] limiter_002_cmd_src_data;                                                                           // limiter_002:cmd_src_data -> cmd_xbar_demux_005:sink_data
	wire   [54:0] limiter_002_cmd_src_channel;                                                                        // limiter_002:cmd_src_channel -> cmd_xbar_demux_005:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                          // cmd_xbar_demux_005:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_mux_005_src_endofpacket;                                                                   // rsp_xbar_mux_005:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_mux_005_src_valid;                                                                         // rsp_xbar_mux_005:src_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_mux_005_src_startofpacket;                                                                 // rsp_xbar_mux_005:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_005_src_data;                                                                          // rsp_xbar_mux_005:src_data -> limiter_002:rsp_sink_data
	wire   [54:0] rsp_xbar_mux_005_src_channel;                                                                       // rsp_xbar_mux_005:src_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_mux_005_src_ready;                                                                         // limiter_002:rsp_sink_ready -> rsp_xbar_mux_005:src_ready
	wire          addr_router_006_src_endofpacket;                                                                    // addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire          addr_router_006_src_valid;                                                                          // addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	wire          addr_router_006_src_startofpacket;                                                                  // addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire  [106:0] addr_router_006_src_data;                                                                           // addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	wire   [54:0] addr_router_006_src_channel;                                                                        // addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	wire          addr_router_006_src_ready;                                                                          // cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	wire          rsp_xbar_mux_006_src_endofpacket;                                                                   // rsp_xbar_mux_006:src_endofpacket -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_006_src_valid;                                                                         // rsp_xbar_mux_006:src_valid -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_006_src_startofpacket;                                                                 // rsp_xbar_mux_006:src_startofpacket -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_006_src_data;                                                                          // rsp_xbar_mux_006:src_data -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] rsp_xbar_mux_006_src_channel;                                                                       // rsp_xbar_mux_006:src_channel -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_006_src_ready;                                                                         // cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_006:src_ready
	wire          addr_router_007_src_endofpacket;                                                                    // addr_router_007:src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	wire          addr_router_007_src_valid;                                                                          // addr_router_007:src_valid -> cmd_xbar_demux_007:sink_valid
	wire          addr_router_007_src_startofpacket;                                                                  // addr_router_007:src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	wire  [106:0] addr_router_007_src_data;                                                                           // addr_router_007:src_data -> cmd_xbar_demux_007:sink_data
	wire   [54:0] addr_router_007_src_channel;                                                                        // addr_router_007:src_channel -> cmd_xbar_demux_007:sink_channel
	wire          addr_router_007_src_ready;                                                                          // cmd_xbar_demux_007:sink_ready -> addr_router_007:src_ready
	wire          rsp_xbar_mux_007_src_endofpacket;                                                                   // rsp_xbar_mux_007:src_endofpacket -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_007_src_valid;                                                                         // rsp_xbar_mux_007:src_valid -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_007_src_startofpacket;                                                                 // rsp_xbar_mux_007:src_startofpacket -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_007_src_data;                                                                          // rsp_xbar_mux_007:src_data -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] rsp_xbar_mux_007_src_channel;                                                                       // rsp_xbar_mux_007:src_channel -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_007_src_ready;                                                                         // cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_007:src_ready
	wire          addr_router_008_src_endofpacket;                                                                    // addr_router_008:src_endofpacket -> cmd_xbar_demux_008:sink_endofpacket
	wire          addr_router_008_src_valid;                                                                          // addr_router_008:src_valid -> cmd_xbar_demux_008:sink_valid
	wire          addr_router_008_src_startofpacket;                                                                  // addr_router_008:src_startofpacket -> cmd_xbar_demux_008:sink_startofpacket
	wire  [106:0] addr_router_008_src_data;                                                                           // addr_router_008:src_data -> cmd_xbar_demux_008:sink_data
	wire   [54:0] addr_router_008_src_channel;                                                                        // addr_router_008:src_channel -> cmd_xbar_demux_008:sink_channel
	wire          addr_router_008_src_ready;                                                                          // cmd_xbar_demux_008:sink_ready -> addr_router_008:src_ready
	wire          rsp_xbar_mux_008_src_endofpacket;                                                                   // rsp_xbar_mux_008:src_endofpacket -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_008_src_valid;                                                                         // rsp_xbar_mux_008:src_valid -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_008_src_startofpacket;                                                                 // rsp_xbar_mux_008:src_startofpacket -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_008_src_data;                                                                          // rsp_xbar_mux_008:src_data -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [54:0] rsp_xbar_mux_008_src_channel;                                                                       // rsp_xbar_mux_008:src_channel -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_008_src_ready;                                                                         // cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_008:src_ready
	wire          limiter_003_cmd_src_endofpacket;                                                                    // limiter_003:cmd_src_endofpacket -> cmd_xbar_demux_009:sink_endofpacket
	wire          limiter_003_cmd_src_startofpacket;                                                                  // limiter_003:cmd_src_startofpacket -> cmd_xbar_demux_009:sink_startofpacket
	wire  [106:0] limiter_003_cmd_src_data;                                                                           // limiter_003:cmd_src_data -> cmd_xbar_demux_009:sink_data
	wire   [54:0] limiter_003_cmd_src_channel;                                                                        // limiter_003:cmd_src_channel -> cmd_xbar_demux_009:sink_channel
	wire          limiter_003_cmd_src_ready;                                                                          // cmd_xbar_demux_009:sink_ready -> limiter_003:cmd_src_ready
	wire          rsp_xbar_mux_009_src_endofpacket;                                                                   // rsp_xbar_mux_009:src_endofpacket -> limiter_003:rsp_sink_endofpacket
	wire          rsp_xbar_mux_009_src_valid;                                                                         // rsp_xbar_mux_009:src_valid -> limiter_003:rsp_sink_valid
	wire          rsp_xbar_mux_009_src_startofpacket;                                                                 // rsp_xbar_mux_009:src_startofpacket -> limiter_003:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_009_src_data;                                                                          // rsp_xbar_mux_009:src_data -> limiter_003:rsp_sink_data
	wire   [54:0] rsp_xbar_mux_009_src_channel;                                                                       // rsp_xbar_mux_009:src_channel -> limiter_003:rsp_sink_channel
	wire          rsp_xbar_mux_009_src_ready;                                                                         // limiter_003:rsp_sink_ready -> rsp_xbar_mux_009:src_ready
	wire          limiter_004_cmd_src_endofpacket;                                                                    // limiter_004:cmd_src_endofpacket -> cmd_xbar_demux_010:sink_endofpacket
	wire          limiter_004_cmd_src_startofpacket;                                                                  // limiter_004:cmd_src_startofpacket -> cmd_xbar_demux_010:sink_startofpacket
	wire  [106:0] limiter_004_cmd_src_data;                                                                           // limiter_004:cmd_src_data -> cmd_xbar_demux_010:sink_data
	wire   [54:0] limiter_004_cmd_src_channel;                                                                        // limiter_004:cmd_src_channel -> cmd_xbar_demux_010:sink_channel
	wire          limiter_004_cmd_src_ready;                                                                          // cmd_xbar_demux_010:sink_ready -> limiter_004:cmd_src_ready
	wire          rsp_xbar_mux_010_src_endofpacket;                                                                   // rsp_xbar_mux_010:src_endofpacket -> limiter_004:rsp_sink_endofpacket
	wire          rsp_xbar_mux_010_src_valid;                                                                         // rsp_xbar_mux_010:src_valid -> limiter_004:rsp_sink_valid
	wire          rsp_xbar_mux_010_src_startofpacket;                                                                 // rsp_xbar_mux_010:src_startofpacket -> limiter_004:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_010_src_data;                                                                          // rsp_xbar_mux_010:src_data -> limiter_004:rsp_sink_data
	wire   [54:0] rsp_xbar_mux_010_src_channel;                                                                       // rsp_xbar_mux_010:src_channel -> limiter_004:rsp_sink_channel
	wire          rsp_xbar_mux_010_src_ready;                                                                         // limiter_004:rsp_sink_ready -> rsp_xbar_mux_010:src_ready
	wire          limiter_005_cmd_src_endofpacket;                                                                    // limiter_005:cmd_src_endofpacket -> cmd_xbar_demux_011:sink_endofpacket
	wire          limiter_005_cmd_src_startofpacket;                                                                  // limiter_005:cmd_src_startofpacket -> cmd_xbar_demux_011:sink_startofpacket
	wire  [106:0] limiter_005_cmd_src_data;                                                                           // limiter_005:cmd_src_data -> cmd_xbar_demux_011:sink_data
	wire   [54:0] limiter_005_cmd_src_channel;                                                                        // limiter_005:cmd_src_channel -> cmd_xbar_demux_011:sink_channel
	wire          limiter_005_cmd_src_ready;                                                                          // cmd_xbar_demux_011:sink_ready -> limiter_005:cmd_src_ready
	wire          rsp_xbar_mux_011_src_endofpacket;                                                                   // rsp_xbar_mux_011:src_endofpacket -> limiter_005:rsp_sink_endofpacket
	wire          rsp_xbar_mux_011_src_valid;                                                                         // rsp_xbar_mux_011:src_valid -> limiter_005:rsp_sink_valid
	wire          rsp_xbar_mux_011_src_startofpacket;                                                                 // rsp_xbar_mux_011:src_startofpacket -> limiter_005:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_011_src_data;                                                                          // rsp_xbar_mux_011:src_data -> limiter_005:rsp_sink_data
	wire   [54:0] rsp_xbar_mux_011_src_channel;                                                                       // rsp_xbar_mux_011:src_channel -> limiter_005:rsp_sink_channel
	wire          rsp_xbar_mux_011_src_ready;                                                                         // limiter_005:rsp_sink_ready -> rsp_xbar_mux_011:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                       // cmd_xbar_mux:src_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                             // cmd_xbar_mux:src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                     // cmd_xbar_mux:src_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_src_data;                                                                              // cmd_xbar_mux:src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_src_channel;                                                                           // cmd_xbar_mux:src_channel -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                          // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                        // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [106:0] id_router_src_data;                                                                                 // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [54:0] id_router_src_channel;                                                                              // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                   // cmd_xbar_mux_001:src_endofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                         // cmd_xbar_mux_001:src_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                 // cmd_xbar_mux_001:src_startofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_001_src_data;                                                                          // cmd_xbar_mux_001:src_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_001_src_channel;                                                                       // cmd_xbar_mux_001:src_channel -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                         // sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                      // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                            // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                    // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [106:0] id_router_001_src_data;                                                                             // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [54:0] id_router_001_src_channel;                                                                          // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_001_src2_ready;                                                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire          id_router_002_src_endofpacket;                                                                      // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                            // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                    // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [106:0] id_router_002_src_data;                                                                             // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [54:0] id_router_002_src_channel;                                                                          // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_003_src_endofpacket;                                                                      // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                            // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                    // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [106:0] id_router_003_src_data;                                                                             // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [54:0] id_router_003_src_channel;                                                                          // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                      // fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                      // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                            // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                    // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [106:0] id_router_004_src_data;                                                                             // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [54:0] id_router_004_src_channel;                                                                          // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                   // cmd_xbar_mux_005:src_endofpacket -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                         // cmd_xbar_mux_005:src_valid -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                 // cmd_xbar_mux_005:src_startofpacket -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_005_src_data;                                                                          // cmd_xbar_mux_005:src_data -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_005_src_channel;                                                                       // cmd_xbar_mux_005:src_channel -> fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                         // fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire          id_router_005_src_endofpacket;                                                                      // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                            // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                    // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [106:0] id_router_005_src_data;                                                                             // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [54:0] id_router_005_src_channel;                                                                          // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                            // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                      // fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                      // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                            // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                    // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [106:0] id_router_006_src_data;                                                                             // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [54:0] id_router_006_src_channel;                                                                          // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                            // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                      // fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                      // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                            // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                    // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [106:0] id_router_007_src_data;                                                                             // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [54:0] id_router_007_src_channel;                                                                          // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                            // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_mux_008_src_endofpacket;                                                                   // cmd_xbar_mux_008:src_endofpacket -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_008_src_valid;                                                                         // cmd_xbar_mux_008:src_valid -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_008_src_startofpacket;                                                                 // cmd_xbar_mux_008:src_startofpacket -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_008_src_data;                                                                          // cmd_xbar_mux_008:src_data -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_008_src_channel;                                                                       // cmd_xbar_mux_008:src_channel -> fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_008_src_ready;                                                                         // fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire          id_router_008_src_endofpacket;                                                                      // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                            // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                    // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [106:0] id_router_008_src_data;                                                                             // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [54:0] id_router_008_src_channel;                                                                          // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                            // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_mux_009_src_endofpacket;                                                                   // cmd_xbar_mux_009:src_endofpacket -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_009_src_valid;                                                                         // cmd_xbar_mux_009:src_valid -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_009_src_startofpacket;                                                                 // cmd_xbar_mux_009:src_startofpacket -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_009_src_data;                                                                          // cmd_xbar_mux_009:src_data -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_009_src_channel;                                                                       // cmd_xbar_mux_009:src_channel -> fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_009_src_ready;                                                                         // fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire          id_router_009_src_endofpacket;                                                                      // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                            // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                    // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [106:0] id_router_009_src_data;                                                                             // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [54:0] id_router_009_src_channel;                                                                          // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                            // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                     // fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_010_src_endofpacket;                                                                      // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                            // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                    // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [106:0] id_router_010_src_data;                                                                             // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [54:0] id_router_010_src_channel;                                                                          // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                            // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_mux_011_src_endofpacket;                                                                   // cmd_xbar_mux_011:src_endofpacket -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_011_src_valid;                                                                         // cmd_xbar_mux_011:src_valid -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_011_src_startofpacket;                                                                 // cmd_xbar_mux_011:src_startofpacket -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_011_src_data;                                                                          // cmd_xbar_mux_011:src_data -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_011_src_channel;                                                                       // cmd_xbar_mux_011:src_channel -> fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_011_src_ready;                                                                         // fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_011:src_ready
	wire          id_router_011_src_endofpacket;                                                                      // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                            // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                    // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [106:0] id_router_011_src_data;                                                                             // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [54:0] id_router_011_src_channel;                                                                          // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                            // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                     // fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                      // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                            // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                    // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [106:0] id_router_012_src_data;                                                                             // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [54:0] id_router_012_src_channel;                                                                          // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                            // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_mux_013_src_endofpacket;                                                                   // cmd_xbar_mux_013:src_endofpacket -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_013_src_valid;                                                                         // cmd_xbar_mux_013:src_valid -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_013_src_startofpacket;                                                                 // cmd_xbar_mux_013:src_startofpacket -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_013_src_data;                                                                          // cmd_xbar_mux_013:src_data -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_013_src_channel;                                                                       // cmd_xbar_mux_013:src_channel -> fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_013_src_ready;                                                                         // fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	wire          id_router_013_src_endofpacket;                                                                      // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                            // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                    // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [106:0] id_router_013_src_data;                                                                             // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [54:0] id_router_013_src_channel;                                                                          // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                            // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_mux_015_src_endofpacket;                                                                   // cmd_xbar_mux_015:src_endofpacket -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_015_src_valid;                                                                         // cmd_xbar_mux_015:src_valid -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_015_src_startofpacket;                                                                 // cmd_xbar_mux_015:src_startofpacket -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_015_src_data;                                                                          // cmd_xbar_mux_015:src_data -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_015_src_channel;                                                                       // cmd_xbar_mux_015:src_channel -> fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_015_src_ready;                                                                         // fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_015:src_ready
	wire          id_router_015_src_endofpacket;                                                                      // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                            // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                    // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [106:0] id_router_015_src_data;                                                                             // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [54:0] id_router_015_src_channel;                                                                          // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                            // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_001_src16_ready;                                                                     // pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire          id_router_016_src_endofpacket;                                                                      // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                            // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                    // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [106:0] id_router_016_src_data;                                                                             // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [54:0] id_router_016_src_channel;                                                                          // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                            // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_mux_017_src_endofpacket;                                                                   // cmd_xbar_mux_017:src_endofpacket -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_017_src_valid;                                                                         // cmd_xbar_mux_017:src_valid -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_017_src_startofpacket;                                                                 // cmd_xbar_mux_017:src_startofpacket -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_017_src_data;                                                                          // cmd_xbar_mux_017:src_data -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_017_src_channel;                                                                       // cmd_xbar_mux_017:src_channel -> instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_017_src_ready;                                                                         // instruction_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_017:src_ready
	wire          id_router_017_src_endofpacket;                                                                      // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                            // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                    // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [106:0] id_router_017_src_data;                                                                             // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [54:0] id_router_017_src_channel;                                                                          // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                            // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_mux_018_src_endofpacket;                                                                   // cmd_xbar_mux_018:src_endofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_018_src_valid;                                                                         // cmd_xbar_mux_018:src_valid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_018_src_startofpacket;                                                                 // cmd_xbar_mux_018:src_startofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_018_src_data;                                                                          // cmd_xbar_mux_018:src_data -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_018_src_channel;                                                                       // cmd_xbar_mux_018:src_channel -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_018_src_ready;                                                                         // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_018:src_ready
	wire          id_router_018_src_endofpacket;                                                                      // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                            // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                    // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [106:0] id_router_018_src_data;                                                                             // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [54:0] id_router_018_src_channel;                                                                          // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                            // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_002_src4_ready;                                                                      // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src4_ready
	wire          id_router_019_src_endofpacket;                                                                      // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                            // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                    // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [106:0] id_router_019_src_data;                                                                             // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [54:0] id_router_019_src_channel;                                                                          // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                            // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          cmd_xbar_demux_002_src5_ready;                                                                      // timer_5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src5_ready
	wire          id_router_020_src_endofpacket;                                                                      // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                            // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                    // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [106:0] id_router_020_src_data;                                                                             // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [54:0] id_router_020_src_channel;                                                                          // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                            // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_demux_002_src7_ready;                                                                      // fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src7_ready
	wire          id_router_022_src_endofpacket;                                                                      // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                            // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                    // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [106:0] id_router_022_src_data;                                                                             // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [54:0] id_router_022_src_channel;                                                                          // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                            // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          cmd_xbar_mux_023_src_endofpacket;                                                                   // cmd_xbar_mux_023:src_endofpacket -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_023_src_valid;                                                                         // cmd_xbar_mux_023:src_valid -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_023_src_startofpacket;                                                                 // cmd_xbar_mux_023:src_startofpacket -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_023_src_data;                                                                          // cmd_xbar_mux_023:src_data -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_023_src_channel;                                                                       // cmd_xbar_mux_023:src_channel -> fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_023_src_ready;                                                                         // fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_023:src_ready
	wire          id_router_023_src_endofpacket;                                                                      // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire          id_router_023_src_valid;                                                                            // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire          id_router_023_src_startofpacket;                                                                    // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [106:0] id_router_023_src_data;                                                                             // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire   [54:0] id_router_023_src_channel;                                                                          // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire          id_router_023_src_ready;                                                                            // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire          cmd_xbar_mux_024_src_endofpacket;                                                                   // cmd_xbar_mux_024:src_endofpacket -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_024_src_valid;                                                                         // cmd_xbar_mux_024:src_valid -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_024_src_startofpacket;                                                                 // cmd_xbar_mux_024:src_startofpacket -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_024_src_data;                                                                          // cmd_xbar_mux_024:src_data -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_024_src_channel;                                                                       // cmd_xbar_mux_024:src_channel -> fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_024_src_ready;                                                                         // fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_024:src_ready
	wire          id_router_024_src_endofpacket;                                                                      // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire          id_router_024_src_valid;                                                                            // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire          id_router_024_src_startofpacket;                                                                    // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [106:0] id_router_024_src_data;                                                                             // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire   [54:0] id_router_024_src_channel;                                                                          // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire          id_router_024_src_ready;                                                                            // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire          cmd_xbar_mux_025_src_endofpacket;                                                                   // cmd_xbar_mux_025:src_endofpacket -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_025_src_valid;                                                                         // cmd_xbar_mux_025:src_valid -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_025_src_startofpacket;                                                                 // cmd_xbar_mux_025:src_startofpacket -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_025_src_data;                                                                          // cmd_xbar_mux_025:src_data -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_025_src_channel;                                                                       // cmd_xbar_mux_025:src_channel -> instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_025_src_ready;                                                                         // instruction_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_025:src_ready
	wire          id_router_025_src_endofpacket;                                                                      // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire          id_router_025_src_valid;                                                                            // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire          id_router_025_src_startofpacket;                                                                    // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire  [106:0] id_router_025_src_data;                                                                             // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire   [54:0] id_router_025_src_channel;                                                                          // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire          id_router_025_src_ready;                                                                            // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire          cmd_xbar_mux_026_src_endofpacket;                                                                   // cmd_xbar_mux_026:src_endofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_026_src_valid;                                                                         // cmd_xbar_mux_026:src_valid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_026_src_startofpacket;                                                                 // cmd_xbar_mux_026:src_startofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_026_src_data;                                                                          // cmd_xbar_mux_026:src_data -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_026_src_channel;                                                                       // cmd_xbar_mux_026:src_channel -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_026_src_ready;                                                                         // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_026:src_ready
	wire          id_router_026_src_endofpacket;                                                                      // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire          id_router_026_src_valid;                                                                            // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire          id_router_026_src_startofpacket;                                                                    // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire  [106:0] id_router_026_src_data;                                                                             // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire   [54:0] id_router_026_src_channel;                                                                          // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire          id_router_026_src_ready;                                                                            // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire          cmd_xbar_demux_003_src6_ready;                                                                      // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src6_ready
	wire          id_router_027_src_endofpacket;                                                                      // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire          id_router_027_src_valid;                                                                            // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire          id_router_027_src_startofpacket;                                                                    // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire  [106:0] id_router_027_src_data;                                                                             // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire   [54:0] id_router_027_src_channel;                                                                          // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire          id_router_027_src_ready;                                                                            // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire          cmd_xbar_demux_003_src7_ready;                                                                      // timer_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src7_ready
	wire          id_router_028_src_endofpacket;                                                                      // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire          id_router_028_src_valid;                                                                            // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire          id_router_028_src_startofpacket;                                                                    // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire  [106:0] id_router_028_src_data;                                                                             // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire   [54:0] id_router_028_src_channel;                                                                          // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire          id_router_028_src_ready;                                                                            // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire          cmd_xbar_demux_003_src8_ready;                                                                      // fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src8_ready
	wire          id_router_029_src_endofpacket;                                                                      // id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire          id_router_029_src_valid;                                                                            // id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	wire          id_router_029_src_startofpacket;                                                                    // id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire  [106:0] id_router_029_src_data;                                                                             // id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	wire   [54:0] id_router_029_src_channel;                                                                          // id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	wire          id_router_029_src_ready;                                                                            // rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	wire          cmd_xbar_demux_003_src9_ready;                                                                      // fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src9_ready
	wire          id_router_030_src_endofpacket;                                                                      // id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire          id_router_030_src_valid;                                                                            // id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	wire          id_router_030_src_startofpacket;                                                                    // id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire  [106:0] id_router_030_src_data;                                                                             // id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	wire   [54:0] id_router_030_src_channel;                                                                          // id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	wire          id_router_030_src_ready;                                                                            // rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	wire          cmd_xbar_demux_003_src10_ready;                                                                     // fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src10_ready
	wire          id_router_031_src_endofpacket;                                                                      // id_router_031:src_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	wire          id_router_031_src_valid;                                                                            // id_router_031:src_valid -> rsp_xbar_demux_031:sink_valid
	wire          id_router_031_src_startofpacket;                                                                    // id_router_031:src_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	wire  [106:0] id_router_031_src_data;                                                                             // id_router_031:src_data -> rsp_xbar_demux_031:sink_data
	wire   [54:0] id_router_031_src_channel;                                                                          // id_router_031:src_channel -> rsp_xbar_demux_031:sink_channel
	wire          id_router_031_src_ready;                                                                            // rsp_xbar_demux_031:sink_ready -> id_router_031:src_ready
	wire          cmd_xbar_mux_032_src_endofpacket;                                                                   // cmd_xbar_mux_032:src_endofpacket -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_032_src_valid;                                                                         // cmd_xbar_mux_032:src_valid -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_032_src_startofpacket;                                                                 // cmd_xbar_mux_032:src_startofpacket -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_032_src_data;                                                                          // cmd_xbar_mux_032:src_data -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_032_src_channel;                                                                       // cmd_xbar_mux_032:src_channel -> instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_032_src_ready;                                                                         // instruction_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_032:src_ready
	wire          id_router_032_src_endofpacket;                                                                      // id_router_032:src_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	wire          id_router_032_src_valid;                                                                            // id_router_032:src_valid -> rsp_xbar_demux_032:sink_valid
	wire          id_router_032_src_startofpacket;                                                                    // id_router_032:src_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	wire  [106:0] id_router_032_src_data;                                                                             // id_router_032:src_data -> rsp_xbar_demux_032:sink_data
	wire   [54:0] id_router_032_src_channel;                                                                          // id_router_032:src_channel -> rsp_xbar_demux_032:sink_channel
	wire          id_router_032_src_ready;                                                                            // rsp_xbar_demux_032:sink_ready -> id_router_032:src_ready
	wire          cmd_xbar_mux_033_src_endofpacket;                                                                   // cmd_xbar_mux_033:src_endofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_033_src_valid;                                                                         // cmd_xbar_mux_033:src_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_033_src_startofpacket;                                                                 // cmd_xbar_mux_033:src_startofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_033_src_data;                                                                          // cmd_xbar_mux_033:src_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_033_src_channel;                                                                       // cmd_xbar_mux_033:src_channel -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_033_src_ready;                                                                         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_033:src_ready
	wire          id_router_033_src_endofpacket;                                                                      // id_router_033:src_endofpacket -> rsp_xbar_demux_033:sink_endofpacket
	wire          id_router_033_src_valid;                                                                            // id_router_033:src_valid -> rsp_xbar_demux_033:sink_valid
	wire          id_router_033_src_startofpacket;                                                                    // id_router_033:src_startofpacket -> rsp_xbar_demux_033:sink_startofpacket
	wire  [106:0] id_router_033_src_data;                                                                             // id_router_033:src_data -> rsp_xbar_demux_033:sink_data
	wire   [54:0] id_router_033_src_channel;                                                                          // id_router_033:src_channel -> rsp_xbar_demux_033:sink_channel
	wire          id_router_033_src_ready;                                                                            // rsp_xbar_demux_033:sink_ready -> id_router_033:src_ready
	wire          cmd_xbar_demux_006_src6_ready;                                                                      // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src6_ready
	wire          id_router_034_src_endofpacket;                                                                      // id_router_034:src_endofpacket -> rsp_xbar_demux_034:sink_endofpacket
	wire          id_router_034_src_valid;                                                                            // id_router_034:src_valid -> rsp_xbar_demux_034:sink_valid
	wire          id_router_034_src_startofpacket;                                                                    // id_router_034:src_startofpacket -> rsp_xbar_demux_034:sink_startofpacket
	wire  [106:0] id_router_034_src_data;                                                                             // id_router_034:src_data -> rsp_xbar_demux_034:sink_data
	wire   [54:0] id_router_034_src_channel;                                                                          // id_router_034:src_channel -> rsp_xbar_demux_034:sink_channel
	wire          id_router_034_src_ready;                                                                            // rsp_xbar_demux_034:sink_ready -> id_router_034:src_ready
	wire          cmd_xbar_demux_006_src7_ready;                                                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src7_ready
	wire          id_router_035_src_endofpacket;                                                                      // id_router_035:src_endofpacket -> rsp_xbar_demux_035:sink_endofpacket
	wire          id_router_035_src_valid;                                                                            // id_router_035:src_valid -> rsp_xbar_demux_035:sink_valid
	wire          id_router_035_src_startofpacket;                                                                    // id_router_035:src_startofpacket -> rsp_xbar_demux_035:sink_startofpacket
	wire  [106:0] id_router_035_src_data;                                                                             // id_router_035:src_data -> rsp_xbar_demux_035:sink_data
	wire   [54:0] id_router_035_src_channel;                                                                          // id_router_035:src_channel -> rsp_xbar_demux_035:sink_channel
	wire          id_router_035_src_ready;                                                                            // rsp_xbar_demux_035:sink_ready -> id_router_035:src_ready
	wire          cmd_xbar_demux_006_src8_ready;                                                                      // fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src8_ready
	wire          id_router_036_src_endofpacket;                                                                      // id_router_036:src_endofpacket -> rsp_xbar_demux_036:sink_endofpacket
	wire          id_router_036_src_valid;                                                                            // id_router_036:src_valid -> rsp_xbar_demux_036:sink_valid
	wire          id_router_036_src_startofpacket;                                                                    // id_router_036:src_startofpacket -> rsp_xbar_demux_036:sink_startofpacket
	wire  [106:0] id_router_036_src_data;                                                                             // id_router_036:src_data -> rsp_xbar_demux_036:sink_data
	wire   [54:0] id_router_036_src_channel;                                                                          // id_router_036:src_channel -> rsp_xbar_demux_036:sink_channel
	wire          id_router_036_src_ready;                                                                            // rsp_xbar_demux_036:sink_ready -> id_router_036:src_ready
	wire          cmd_xbar_demux_006_src9_ready;                                                                      // fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src9_ready
	wire          id_router_037_src_endofpacket;                                                                      // id_router_037:src_endofpacket -> rsp_xbar_demux_037:sink_endofpacket
	wire          id_router_037_src_valid;                                                                            // id_router_037:src_valid -> rsp_xbar_demux_037:sink_valid
	wire          id_router_037_src_startofpacket;                                                                    // id_router_037:src_startofpacket -> rsp_xbar_demux_037:sink_startofpacket
	wire  [106:0] id_router_037_src_data;                                                                             // id_router_037:src_data -> rsp_xbar_demux_037:sink_data
	wire   [54:0] id_router_037_src_channel;                                                                          // id_router_037:src_channel -> rsp_xbar_demux_037:sink_channel
	wire          id_router_037_src_ready;                                                                            // rsp_xbar_demux_037:sink_ready -> id_router_037:src_ready
	wire          cmd_xbar_demux_006_src10_ready;                                                                     // fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src10_ready
	wire          id_router_038_src_endofpacket;                                                                      // id_router_038:src_endofpacket -> rsp_xbar_demux_038:sink_endofpacket
	wire          id_router_038_src_valid;                                                                            // id_router_038:src_valid -> rsp_xbar_demux_038:sink_valid
	wire          id_router_038_src_startofpacket;                                                                    // id_router_038:src_startofpacket -> rsp_xbar_demux_038:sink_startofpacket
	wire  [106:0] id_router_038_src_data;                                                                             // id_router_038:src_data -> rsp_xbar_demux_038:sink_data
	wire   [54:0] id_router_038_src_channel;                                                                          // id_router_038:src_channel -> rsp_xbar_demux_038:sink_channel
	wire          id_router_038_src_ready;                                                                            // rsp_xbar_demux_038:sink_ready -> id_router_038:src_ready
	wire          cmd_xbar_demux_006_src11_ready;                                                                     // fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src11_ready
	wire          id_router_039_src_endofpacket;                                                                      // id_router_039:src_endofpacket -> rsp_xbar_demux_039:sink_endofpacket
	wire          id_router_039_src_valid;                                                                            // id_router_039:src_valid -> rsp_xbar_demux_039:sink_valid
	wire          id_router_039_src_startofpacket;                                                                    // id_router_039:src_startofpacket -> rsp_xbar_demux_039:sink_startofpacket
	wire  [106:0] id_router_039_src_data;                                                                             // id_router_039:src_data -> rsp_xbar_demux_039:sink_data
	wire   [54:0] id_router_039_src_channel;                                                                          // id_router_039:src_channel -> rsp_xbar_demux_039:sink_channel
	wire          id_router_039_src_ready;                                                                            // rsp_xbar_demux_039:sink_ready -> id_router_039:src_ready
	wire          cmd_xbar_mux_040_src_endofpacket;                                                                   // cmd_xbar_mux_040:src_endofpacket -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_040_src_valid;                                                                         // cmd_xbar_mux_040:src_valid -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_040_src_startofpacket;                                                                 // cmd_xbar_mux_040:src_startofpacket -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_040_src_data;                                                                          // cmd_xbar_mux_040:src_data -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_040_src_channel;                                                                       // cmd_xbar_mux_040:src_channel -> fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_040_src_ready;                                                                         // fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_040:src_ready
	wire          id_router_040_src_endofpacket;                                                                      // id_router_040:src_endofpacket -> rsp_xbar_demux_040:sink_endofpacket
	wire          id_router_040_src_valid;                                                                            // id_router_040:src_valid -> rsp_xbar_demux_040:sink_valid
	wire          id_router_040_src_startofpacket;                                                                    // id_router_040:src_startofpacket -> rsp_xbar_demux_040:sink_startofpacket
	wire  [106:0] id_router_040_src_data;                                                                             // id_router_040:src_data -> rsp_xbar_demux_040:sink_data
	wire   [54:0] id_router_040_src_channel;                                                                          // id_router_040:src_channel -> rsp_xbar_demux_040:sink_channel
	wire          id_router_040_src_ready;                                                                            // rsp_xbar_demux_040:sink_ready -> id_router_040:src_ready
	wire          cmd_xbar_mux_041_src_endofpacket;                                                                   // cmd_xbar_mux_041:src_endofpacket -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_041_src_valid;                                                                         // cmd_xbar_mux_041:src_valid -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_041_src_startofpacket;                                                                 // cmd_xbar_mux_041:src_startofpacket -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_041_src_data;                                                                          // cmd_xbar_mux_041:src_data -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_041_src_channel;                                                                       // cmd_xbar_mux_041:src_channel -> instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_041_src_ready;                                                                         // instruction_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_041:src_ready
	wire          id_router_041_src_endofpacket;                                                                      // id_router_041:src_endofpacket -> rsp_xbar_demux_041:sink_endofpacket
	wire          id_router_041_src_valid;                                                                            // id_router_041:src_valid -> rsp_xbar_demux_041:sink_valid
	wire          id_router_041_src_startofpacket;                                                                    // id_router_041:src_startofpacket -> rsp_xbar_demux_041:sink_startofpacket
	wire  [106:0] id_router_041_src_data;                                                                             // id_router_041:src_data -> rsp_xbar_demux_041:sink_data
	wire   [54:0] id_router_041_src_channel;                                                                          // id_router_041:src_channel -> rsp_xbar_demux_041:sink_channel
	wire          id_router_041_src_ready;                                                                            // rsp_xbar_demux_041:sink_ready -> id_router_041:src_ready
	wire          cmd_xbar_mux_042_src_endofpacket;                                                                   // cmd_xbar_mux_042:src_endofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_042_src_valid;                                                                         // cmd_xbar_mux_042:src_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_042_src_startofpacket;                                                                 // cmd_xbar_mux_042:src_startofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_042_src_data;                                                                          // cmd_xbar_mux_042:src_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_042_src_channel;                                                                       // cmd_xbar_mux_042:src_channel -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_042_src_ready;                                                                         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_042:src_ready
	wire          id_router_042_src_endofpacket;                                                                      // id_router_042:src_endofpacket -> rsp_xbar_demux_042:sink_endofpacket
	wire          id_router_042_src_valid;                                                                            // id_router_042:src_valid -> rsp_xbar_demux_042:sink_valid
	wire          id_router_042_src_startofpacket;                                                                    // id_router_042:src_startofpacket -> rsp_xbar_demux_042:sink_startofpacket
	wire  [106:0] id_router_042_src_data;                                                                             // id_router_042:src_data -> rsp_xbar_demux_042:sink_data
	wire   [54:0] id_router_042_src_channel;                                                                          // id_router_042:src_channel -> rsp_xbar_demux_042:sink_channel
	wire          id_router_042_src_ready;                                                                            // rsp_xbar_demux_042:sink_ready -> id_router_042:src_ready
	wire          cmd_xbar_demux_007_src4_ready;                                                                      // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src4_ready
	wire          id_router_043_src_endofpacket;                                                                      // id_router_043:src_endofpacket -> rsp_xbar_demux_043:sink_endofpacket
	wire          id_router_043_src_valid;                                                                            // id_router_043:src_valid -> rsp_xbar_demux_043:sink_valid
	wire          id_router_043_src_startofpacket;                                                                    // id_router_043:src_startofpacket -> rsp_xbar_demux_043:sink_startofpacket
	wire  [106:0] id_router_043_src_data;                                                                             // id_router_043:src_data -> rsp_xbar_demux_043:sink_data
	wire   [54:0] id_router_043_src_channel;                                                                          // id_router_043:src_channel -> rsp_xbar_demux_043:sink_channel
	wire          id_router_043_src_ready;                                                                            // rsp_xbar_demux_043:sink_ready -> id_router_043:src_ready
	wire          cmd_xbar_demux_007_src5_ready;                                                                      // timer_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src5_ready
	wire          id_router_044_src_endofpacket;                                                                      // id_router_044:src_endofpacket -> rsp_xbar_demux_044:sink_endofpacket
	wire          id_router_044_src_valid;                                                                            // id_router_044:src_valid -> rsp_xbar_demux_044:sink_valid
	wire          id_router_044_src_startofpacket;                                                                    // id_router_044:src_startofpacket -> rsp_xbar_demux_044:sink_startofpacket
	wire  [106:0] id_router_044_src_data;                                                                             // id_router_044:src_data -> rsp_xbar_demux_044:sink_data
	wire   [54:0] id_router_044_src_channel;                                                                          // id_router_044:src_channel -> rsp_xbar_demux_044:sink_channel
	wire          id_router_044_src_ready;                                                                            // rsp_xbar_demux_044:sink_ready -> id_router_044:src_ready
	wire          cmd_xbar_demux_007_src6_ready;                                                                      // fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src6_ready
	wire          id_router_045_src_endofpacket;                                                                      // id_router_045:src_endofpacket -> rsp_xbar_demux_045:sink_endofpacket
	wire          id_router_045_src_valid;                                                                            // id_router_045:src_valid -> rsp_xbar_demux_045:sink_valid
	wire          id_router_045_src_startofpacket;                                                                    // id_router_045:src_startofpacket -> rsp_xbar_demux_045:sink_startofpacket
	wire  [106:0] id_router_045_src_data;                                                                             // id_router_045:src_data -> rsp_xbar_demux_045:sink_data
	wire   [54:0] id_router_045_src_channel;                                                                          // id_router_045:src_channel -> rsp_xbar_demux_045:sink_channel
	wire          id_router_045_src_ready;                                                                            // rsp_xbar_demux_045:sink_ready -> id_router_045:src_ready
	wire          cmd_xbar_demux_007_src7_ready;                                                                      // fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src7_ready
	wire          id_router_046_src_endofpacket;                                                                      // id_router_046:src_endofpacket -> rsp_xbar_demux_046:sink_endofpacket
	wire          id_router_046_src_valid;                                                                            // id_router_046:src_valid -> rsp_xbar_demux_046:sink_valid
	wire          id_router_046_src_startofpacket;                                                                    // id_router_046:src_startofpacket -> rsp_xbar_demux_046:sink_startofpacket
	wire  [106:0] id_router_046_src_data;                                                                             // id_router_046:src_data -> rsp_xbar_demux_046:sink_data
	wire   [54:0] id_router_046_src_channel;                                                                          // id_router_046:src_channel -> rsp_xbar_demux_046:sink_channel
	wire          id_router_046_src_ready;                                                                            // rsp_xbar_demux_046:sink_ready -> id_router_046:src_ready
	wire          cmd_xbar_mux_047_src_endofpacket;                                                                   // cmd_xbar_mux_047:src_endofpacket -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_047_src_valid;                                                                         // cmd_xbar_mux_047:src_valid -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_047_src_startofpacket;                                                                 // cmd_xbar_mux_047:src_startofpacket -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_047_src_data;                                                                          // cmd_xbar_mux_047:src_data -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_047_src_channel;                                                                       // cmd_xbar_mux_047:src_channel -> fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_047_src_ready;                                                                         // fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_047:src_ready
	wire          id_router_047_src_endofpacket;                                                                      // id_router_047:src_endofpacket -> rsp_xbar_demux_047:sink_endofpacket
	wire          id_router_047_src_valid;                                                                            // id_router_047:src_valid -> rsp_xbar_demux_047:sink_valid
	wire          id_router_047_src_startofpacket;                                                                    // id_router_047:src_startofpacket -> rsp_xbar_demux_047:sink_startofpacket
	wire  [106:0] id_router_047_src_data;                                                                             // id_router_047:src_data -> rsp_xbar_demux_047:sink_data
	wire   [54:0] id_router_047_src_channel;                                                                          // id_router_047:src_channel -> rsp_xbar_demux_047:sink_channel
	wire          id_router_047_src_ready;                                                                            // rsp_xbar_demux_047:sink_ready -> id_router_047:src_ready
	wire          cmd_xbar_mux_048_src_endofpacket;                                                                   // cmd_xbar_mux_048:src_endofpacket -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_048_src_valid;                                                                         // cmd_xbar_mux_048:src_valid -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_048_src_startofpacket;                                                                 // cmd_xbar_mux_048:src_startofpacket -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_048_src_data;                                                                          // cmd_xbar_mux_048:src_data -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_048_src_channel;                                                                       // cmd_xbar_mux_048:src_channel -> instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_048_src_ready;                                                                         // instruction_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_048:src_ready
	wire          id_router_048_src_endofpacket;                                                                      // id_router_048:src_endofpacket -> rsp_xbar_demux_048:sink_endofpacket
	wire          id_router_048_src_valid;                                                                            // id_router_048:src_valid -> rsp_xbar_demux_048:sink_valid
	wire          id_router_048_src_startofpacket;                                                                    // id_router_048:src_startofpacket -> rsp_xbar_demux_048:sink_startofpacket
	wire  [106:0] id_router_048_src_data;                                                                             // id_router_048:src_data -> rsp_xbar_demux_048:sink_data
	wire   [54:0] id_router_048_src_channel;                                                                          // id_router_048:src_channel -> rsp_xbar_demux_048:sink_channel
	wire          id_router_048_src_ready;                                                                            // rsp_xbar_demux_048:sink_ready -> id_router_048:src_ready
	wire          cmd_xbar_mux_049_src_endofpacket;                                                                   // cmd_xbar_mux_049:src_endofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_049_src_valid;                                                                         // cmd_xbar_mux_049:src_valid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_049_src_startofpacket;                                                                 // cmd_xbar_mux_049:src_startofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_049_src_data;                                                                          // cmd_xbar_mux_049:src_data -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [54:0] cmd_xbar_mux_049_src_channel;                                                                       // cmd_xbar_mux_049:src_channel -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_049_src_ready;                                                                         // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_049:src_ready
	wire          id_router_049_src_endofpacket;                                                                      // id_router_049:src_endofpacket -> rsp_xbar_demux_049:sink_endofpacket
	wire          id_router_049_src_valid;                                                                            // id_router_049:src_valid -> rsp_xbar_demux_049:sink_valid
	wire          id_router_049_src_startofpacket;                                                                    // id_router_049:src_startofpacket -> rsp_xbar_demux_049:sink_startofpacket
	wire  [106:0] id_router_049_src_data;                                                                             // id_router_049:src_data -> rsp_xbar_demux_049:sink_data
	wire   [54:0] id_router_049_src_channel;                                                                          // id_router_049:src_channel -> rsp_xbar_demux_049:sink_channel
	wire          id_router_049_src_ready;                                                                            // rsp_xbar_demux_049:sink_ready -> id_router_049:src_ready
	wire          cmd_xbar_demux_008_src6_ready;                                                                      // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src6_ready
	wire          id_router_050_src_endofpacket;                                                                      // id_router_050:src_endofpacket -> rsp_xbar_demux_050:sink_endofpacket
	wire          id_router_050_src_valid;                                                                            // id_router_050:src_valid -> rsp_xbar_demux_050:sink_valid
	wire          id_router_050_src_startofpacket;                                                                    // id_router_050:src_startofpacket -> rsp_xbar_demux_050:sink_startofpacket
	wire  [106:0] id_router_050_src_data;                                                                             // id_router_050:src_data -> rsp_xbar_demux_050:sink_data
	wire   [54:0] id_router_050_src_channel;                                                                          // id_router_050:src_channel -> rsp_xbar_demux_050:sink_channel
	wire          id_router_050_src_ready;                                                                            // rsp_xbar_demux_050:sink_ready -> id_router_050:src_ready
	wire          cmd_xbar_demux_008_src7_ready;                                                                      // timer_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src7_ready
	wire          id_router_051_src_endofpacket;                                                                      // id_router_051:src_endofpacket -> rsp_xbar_demux_051:sink_endofpacket
	wire          id_router_051_src_valid;                                                                            // id_router_051:src_valid -> rsp_xbar_demux_051:sink_valid
	wire          id_router_051_src_startofpacket;                                                                    // id_router_051:src_startofpacket -> rsp_xbar_demux_051:sink_startofpacket
	wire  [106:0] id_router_051_src_data;                                                                             // id_router_051:src_data -> rsp_xbar_demux_051:sink_data
	wire   [54:0] id_router_051_src_channel;                                                                          // id_router_051:src_channel -> rsp_xbar_demux_051:sink_channel
	wire          id_router_051_src_ready;                                                                            // rsp_xbar_demux_051:sink_ready -> id_router_051:src_ready
	wire          cmd_xbar_demux_008_src8_ready;                                                                      // fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src8_ready
	wire          id_router_052_src_endofpacket;                                                                      // id_router_052:src_endofpacket -> rsp_xbar_demux_052:sink_endofpacket
	wire          id_router_052_src_valid;                                                                            // id_router_052:src_valid -> rsp_xbar_demux_052:sink_valid
	wire          id_router_052_src_startofpacket;                                                                    // id_router_052:src_startofpacket -> rsp_xbar_demux_052:sink_startofpacket
	wire  [106:0] id_router_052_src_data;                                                                             // id_router_052:src_data -> rsp_xbar_demux_052:sink_data
	wire   [54:0] id_router_052_src_channel;                                                                          // id_router_052:src_channel -> rsp_xbar_demux_052:sink_channel
	wire          id_router_052_src_ready;                                                                            // rsp_xbar_demux_052:sink_ready -> id_router_052:src_ready
	wire          cmd_xbar_demux_008_src9_ready;                                                                      // fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src9_ready
	wire          id_router_053_src_endofpacket;                                                                      // id_router_053:src_endofpacket -> rsp_xbar_demux_053:sink_endofpacket
	wire          id_router_053_src_valid;                                                                            // id_router_053:src_valid -> rsp_xbar_demux_053:sink_valid
	wire          id_router_053_src_startofpacket;                                                                    // id_router_053:src_startofpacket -> rsp_xbar_demux_053:sink_startofpacket
	wire  [106:0] id_router_053_src_data;                                                                             // id_router_053:src_data -> rsp_xbar_demux_053:sink_data
	wire   [54:0] id_router_053_src_channel;                                                                          // id_router_053:src_channel -> rsp_xbar_demux_053:sink_channel
	wire          id_router_053_src_ready;                                                                            // rsp_xbar_demux_053:sink_ready -> id_router_053:src_ready
	wire          cmd_xbar_demux_008_src10_ready;                                                                     // fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src10_ready
	wire          id_router_054_src_endofpacket;                                                                      // id_router_054:src_endofpacket -> rsp_xbar_demux_054:sink_endofpacket
	wire          id_router_054_src_valid;                                                                            // id_router_054:src_valid -> rsp_xbar_demux_054:sink_valid
	wire          id_router_054_src_startofpacket;                                                                    // id_router_054:src_startofpacket -> rsp_xbar_demux_054:sink_startofpacket
	wire  [106:0] id_router_054_src_data;                                                                             // id_router_054:src_data -> rsp_xbar_demux_054:sink_data
	wire   [54:0] id_router_054_src_channel;                                                                          // id_router_054:src_channel -> rsp_xbar_demux_054:sink_channel
	wire          id_router_054_src_ready;                                                                            // rsp_xbar_demux_054:sink_ready -> id_router_054:src_ready
	wire          cmd_xbar_demux_001_src14_ready;                                                                     // width_adapter:in_ready -> cmd_xbar_demux_001:src14_ready
	wire          width_adapter_src_endofpacket;                                                                      // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                            // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                    // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [79:0] width_adapter_src_data;                                                                             // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                            // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [54:0] width_adapter_src_channel;                                                                          // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_014_src_endofpacket;                                                                      // id_router_014:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_014_src_valid;                                                                            // id_router_014:src_valid -> width_adapter_001:in_valid
	wire          id_router_014_src_startofpacket;                                                                    // id_router_014:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [79:0] id_router_014_src_data;                                                                             // id_router_014:src_data -> width_adapter_001:in_data
	wire   [54:0] id_router_014_src_channel;                                                                          // id_router_014:src_channel -> width_adapter_001:in_channel
	wire          id_router_014_src_ready;                                                                            // width_adapter_001:in_ready -> id_router_014:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                  // width_adapter_001:out_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                        // width_adapter_001:out_valid -> rsp_xbar_demux_014:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                // width_adapter_001:out_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [106:0] width_adapter_001_src_data;                                                                         // width_adapter_001:out_data -> rsp_xbar_demux_014:sink_data
	wire          width_adapter_001_src_ready;                                                                        // rsp_xbar_demux_014:sink_ready -> width_adapter_001:out_ready
	wire   [54:0] width_adapter_001_src_channel;                                                                      // width_adapter_001:out_channel -> rsp_xbar_demux_014:sink_channel
	wire          cmd_xbar_demux_002_src6_ready;                                                                      // width_adapter_002:in_ready -> cmd_xbar_demux_002:src6_ready
	wire          width_adapter_002_src_endofpacket;                                                                  // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                        // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [79:0] width_adapter_002_src_data;                                                                         // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_002_src_ready;                                                                        // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire   [54:0] width_adapter_002_src_channel;                                                                      // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_021_src_endofpacket;                                                                      // id_router_021:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_021_src_valid;                                                                            // id_router_021:src_valid -> width_adapter_003:in_valid
	wire          id_router_021_src_startofpacket;                                                                    // id_router_021:src_startofpacket -> width_adapter_003:in_startofpacket
	wire   [79:0] id_router_021_src_data;                                                                             // id_router_021:src_data -> width_adapter_003:in_data
	wire   [54:0] id_router_021_src_channel;                                                                          // id_router_021:src_channel -> width_adapter_003:in_channel
	wire          id_router_021_src_ready;                                                                            // width_adapter_003:in_ready -> id_router_021:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                  // width_adapter_003:out_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                        // width_adapter_003:out_valid -> rsp_xbar_demux_021:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                                // width_adapter_003:out_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [106:0] width_adapter_003_src_data;                                                                         // width_adapter_003:out_data -> rsp_xbar_demux_021:sink_data
	wire          width_adapter_003_src_ready;                                                                        // rsp_xbar_demux_021:sink_ready -> width_adapter_003:out_ready
	wire   [54:0] width_adapter_003_src_channel;                                                                      // width_adapter_003:out_channel -> rsp_xbar_demux_021:sink_channel
	wire   [54:0] limiter_cmd_valid_data;                                                                             // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [54:0] limiter_001_cmd_valid_data;                                                                         // limiter_001:cmd_src_valid -> cmd_xbar_demux_004:sink_valid
	wire   [54:0] limiter_002_cmd_valid_data;                                                                         // limiter_002:cmd_src_valid -> cmd_xbar_demux_005:sink_valid
	wire   [54:0] limiter_003_cmd_valid_data;                                                                         // limiter_003:cmd_src_valid -> cmd_xbar_demux_009:sink_valid
	wire   [54:0] limiter_004_cmd_valid_data;                                                                         // limiter_004:cmd_src_valid -> cmd_xbar_demux_010:sink_valid
	wire   [54:0] limiter_005_cmd_valid_data;                                                                         // limiter_005:cmd_src_valid -> cmd_xbar_demux_011:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                           // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                           // timer_0:irq -> irq_mapper:receiver1_irq
	wire   [31:0] cpu_0_d_irq_irq;                                                                                    // irq_mapper:sender_irq -> cpu_0:d_irq
	wire          irq_mapper_001_receiver0_irq;                                                                       // jtag_uart_1:av_irq -> irq_mapper_001:receiver0_irq
	wire          irq_mapper_001_receiver1_irq;                                                                       // timer_1:irq -> irq_mapper_001:receiver1_irq
	wire   [31:0] cpu_1_d_irq_irq;                                                                                    // irq_mapper_001:sender_irq -> cpu_1:d_irq
	wire          irq_mapper_002_receiver0_irq;                                                                       // timer_2:irq -> irq_mapper_002:receiver0_irq
	wire          irq_mapper_002_receiver1_irq;                                                                       // jtag_uart_2:av_irq -> irq_mapper_002:receiver1_irq
	wire   [31:0] cpu_2_d_irq_irq;                                                                                    // irq_mapper_002:sender_irq -> cpu_2:d_irq
	wire          irq_mapper_003_receiver0_irq;                                                                       // jtag_uart_3:av_irq -> irq_mapper_003:receiver0_irq
	wire          irq_mapper_003_receiver1_irq;                                                                       // timer_3:irq -> irq_mapper_003:receiver1_irq
	wire   [31:0] cpu_3_d_irq_irq;                                                                                    // irq_mapper_003:sender_irq -> cpu_3:d_irq
	wire          irq_mapper_004_receiver0_irq;                                                                       // timer_4:irq -> irq_mapper_004:receiver0_irq
	wire          irq_mapper_004_receiver1_irq;                                                                       // jtag_uart_4:av_irq -> irq_mapper_004:receiver1_irq
	wire   [31:0] cpu_4_d_irq_irq;                                                                                    // irq_mapper_004:sender_irq -> cpu_4:d_irq
	wire          irq_mapper_005_receiver0_irq;                                                                       // jtag_uart_5:av_irq -> irq_mapper_005:receiver0_irq
	wire          irq_mapper_005_receiver1_irq;                                                                       // timer_5:irq -> irq_mapper_005:receiver1_irq
	wire   [31:0] cpu_5_d_irq_irq;                                                                                    // irq_mapper_005:sender_irq -> cpu_5:d_irq

	SoC_cpu_0 cpu_0 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (cpu_0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_0_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_0_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_0_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_0_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	SoC_timer_0 timer_0 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                              //   irq.irq
	);

	SoC_instruction_mem_1 instruction_mem_1 (
		.clk        (clk_clk),                                                        //   clk1.clk
		.address    (instruction_mem_1_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (instruction_mem_1_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (instruction_mem_1_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (instruction_mem_1_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (instruction_mem_1_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (instruction_mem_1_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (instruction_mem_1_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset)                              // reset1.reset
	);

	SoC_cpu_1 cpu_1 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (cpu_1_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_1_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_1_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_1_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_1_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_1_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_1_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_1_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_1_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_1_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_1_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_1_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_1_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_1 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver0_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_1 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                  // reset.reset_n
		.address    (timer_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_001_receiver1_irq)                          //   irq.irq
	);

	SoC_instruction_mem_2 instruction_mem_2 (
		.clk        (clk_clk),                                                        //   clk1.clk
		.address    (instruction_mem_2_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (instruction_mem_2_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (instruction_mem_2_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (instruction_mem_2_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (instruction_mem_2_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (instruction_mem_2_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (instruction_mem_2_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset)                              // reset1.reset
	);

	SoC_cpu_2 cpu_2 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (cpu_2_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_2_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_2_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_2_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_2_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_2_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_2_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_2_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_2_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_2_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_2_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_2_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_2_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_2_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_2_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_2 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~cpu_2_jtag_debug_module_reset_reset),                                     //             reset.reset_n
		.av_chipselect  (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver1_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_2 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                  // reset.reset_n
		.address    (timer_2_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_2_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_2_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_2_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_2_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_002_receiver0_irq)                          //   irq.irq
	);

	SoC_instruction_mem_3 instruction_mem_3 (
		.clk        (clk_clk),                                                        //   clk1.clk
		.address    (instruction_mem_3_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (instruction_mem_3_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (instruction_mem_3_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (instruction_mem_3_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (instruction_mem_3_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (instruction_mem_3_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (instruction_mem_3_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_004_reset_out_reset)                              // reset1.reset
	);

	SoC_cpu_3 cpu_3 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (cpu_3_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_3_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_3_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_3_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_3_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_3_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_3_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_3_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_3_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_3_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_3_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_3_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_3_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_3_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_3_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_3 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_004_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_003_receiver0_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_3 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                  // reset.reset_n
		.address    (timer_3_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_3_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_3_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_3_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_3_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_003_receiver1_irq)                          //   irq.irq
	);

	SoC_instruction_mem_4 instruction_mem_4 (
		.clk        (clk_clk),                                                        //   clk1.clk
		.address    (instruction_mem_4_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (instruction_mem_4_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (instruction_mem_4_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (instruction_mem_4_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (instruction_mem_4_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (instruction_mem_4_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (instruction_mem_4_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_005_reset_out_reset)                              // reset1.reset
	);

	SoC_cpu_4 cpu_4 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (cpu_4_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_4_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_4_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_4_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_4_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_4_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_4_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_4_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_4_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_4_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_4_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_4_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_4_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_4_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_4_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_4 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_005_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_004_receiver1_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_4 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_005_reset_out_reset),                  // reset.reset_n
		.address    (timer_4_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_4_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_4_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_4_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_4_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_004_receiver0_irq)                          //   irq.irq
	);

	SoC_instruction_mem_5 instruction_mem_5 (
		.clk        (clk_clk),                                                        //   clk1.clk
		.address    (instruction_mem_5_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (instruction_mem_5_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (instruction_mem_5_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (instruction_mem_5_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (instruction_mem_5_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (instruction_mem_5_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (instruction_mem_5_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_006_reset_out_reset)                              // reset1.reset
	);

	SoC_cpu_5 cpu_5 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (cpu_5_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_5_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_5_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_5_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_5_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_5_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_5_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_5_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_5_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_5_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_5_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_5_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_5_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_5_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_5_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_5 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_006_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_005_receiver0_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_5 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),                  // reset.reset_n
		.address    (timer_5_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_5_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_5_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_5_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_5_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_005_receiver1_irq)                          //   irq.irq
	);

	SoC_fifo_0_stage1_to_2 fifo_0_stage1_to_2 (
		.wrclock                          (clk_clk),                                                            //   clk_in.clk
		.reset_n                          (~rst_controller_007_reset_out_reset),                                // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_0_stage1_to_2_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_0_stage1_to_2_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_0_stage1_to_2_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                   //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_0_stage1_to_2_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_0_stage1_to_2_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_0_stage1_to_2_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_fifo_0_stage1_to_2 fifo_1_stage1_to_2 (
		.wrclock                          (clk_clk),                                                            //   clk_in.clk
		.reset_n                          (~rst_controller_007_reset_out_reset),                                // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_1_stage1_to_2_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_1_stage1_to_2_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_1_stage1_to_2_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                   //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_1_stage1_to_2_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_1_stage1_to_2_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_1_stage1_to_2_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_fifo_0_stage1_to_2 fifo_2_stage1_to_2 (
		.wrclock                          (clk_clk),                                                            //   clk_in.clk
		.reset_n                          (~rst_controller_007_reset_out_reset),                                // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_2_stage1_to_2_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_2_stage1_to_2_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_2_stage1_to_2_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                   //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_2_stage1_to_2_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_2_stage1_to_2_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_2_stage1_to_2_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_fifo_stage1_to_4 fifo_stage1_to_4 (
		.wrclock                          (clk_clk),                                                          //   clk_in.clk
		.reset_n                          (~rst_controller_008_reset_out_reset),                              // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_stage1_to_4_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_stage1_to_4_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_stage1_to_4_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                 //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_stage1_to_4_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_stage1_to_4_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_stage1_to_4_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_fifo_stage1_to_4 fifo_stage1_to_5 (
		.wrclock                          (clk_clk),                                                          //   clk_in.clk
		.reset_n                          (~rst_controller_009_reset_out_reset),                              // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_stage1_to_5_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_stage1_to_5_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_stage1_to_5_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                 //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_stage1_to_5_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_stage1_to_5_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_stage1_to_5_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_fifo_stage1_to_6 fifo_stage1_to_6 (
		.wrclock                          (clk_clk),                                                          //   clk_in.clk
		.reset_n                          (~rst_controller_010_reset_out_reset),                              // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_stage1_to_6_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_stage1_to_6_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_stage1_to_6_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                 //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_stage1_to_6_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_stage1_to_6_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_stage1_to_6_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_fifo_stage2_to_3 fifo_stage2_to_3 (
		.wrclock                          (clk_clk),                                                          //   clk_in.clk
		.reset_n                          (~rst_controller_011_reset_out_reset),                              // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_stage2_to_3_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_stage2_to_3_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_stage2_to_3_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                 //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_stage2_to_3_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_stage2_to_3_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_stage2_to_3_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_fifo_stage2_to_3 fifo_stage3_to_4 (
		.wrclock                          (clk_clk),                                                          //   clk_in.clk
		.reset_n                          (~rst_controller_012_reset_out_reset),                              // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_stage3_to_4_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_stage3_to_4_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_stage3_to_4_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                 //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_stage3_to_4_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_stage3_to_4_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_stage3_to_4_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_fifo_stage2_to_3 fifo_stage4_to_5 (
		.wrclock                          (clk_clk),                                                          //   clk_in.clk
		.reset_n                          (~rst_controller_013_reset_out_reset),                              // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_stage4_to_5_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_stage4_to_5_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_stage4_to_5_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                 //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_stage4_to_5_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_stage4_to_5_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_stage4_to_5_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_fifo_stage2_to_3 fifo_stage5_to_6 (
		.wrclock                          (clk_clk),                                                          //   clk_in.clk
		.reset_n                          (~rst_controller_014_reset_out_reset),                              // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_stage5_to_6_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_stage5_to_6_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_stage5_to_6_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (),                                                                 //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_stage5_to_6_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_stage5_to_6_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_stage5_to_6_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_pll pll (
		.clk       (clk_clk),                                                //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),                     // inclk_interface_reset.reset
		.read      (pll_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (pll_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (pll_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (pll_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (pll_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (c0_clk),                                                 //                    c0.clk
		.areset    (),                                                       //        areset_conduit.export
		.locked    (),                                                       //        locked_conduit.export
		.phasedone ()                                                        //     phasedone_conduit.export
	);

	SoC_sdram_controller sdram_controller (
		.clk            (clk_clk),                                                          //   clk.clk
		.reset_n        (~rst_controller_015_reset_out_reset),                              // reset.reset_n
		.az_addr        (sdram_controller_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_controller_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_controller_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_controller_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_controller_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_controller_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_controller_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_controller_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_controller_wire_dq),                                         //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                                        //      .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_0_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_0_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_0_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_0_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_0_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_0_data_master_read),                                               //                          .read
		.av_readdata           (cpu_0_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_0_data_master_write),                                              //                          .write
		.av_writedata          (cpu_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_5_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_5_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_5_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_5_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_5_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_5_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_5_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_5_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_5_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_5_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_5_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_5_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_5_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_5_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_5_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_5_data_master_read),                                               //                          .read
		.av_readdata           (cpu_5_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_5_data_master_write),                                              //                          .write
		.av_writedata          (cpu_5_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_5_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_1_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_1_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_1_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_1_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_1_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_1_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_1_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_1_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_1_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_1_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_1_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_1_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_1_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_1_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_1_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_1_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_1_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_1_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_1_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_1_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_1_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_1_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_1_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_1_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_1_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_1_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_1_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_1_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_1_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_1_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_1_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_1_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_1_data_master_read),                                               //                          .read
		.av_readdata           (cpu_1_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_1_data_master_write),                                              //                          .write
		.av_writedata          (cpu_1_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_1_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_2_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_2_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_2_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_2_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_2_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_2_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_2_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_2_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_2_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_2_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_2_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_2_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_2_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_2_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_2_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_2_data_master_read),                                               //                          .read
		.av_readdata           (cpu_2_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_2_data_master_write),                                              //                          .write
		.av_writedata          (cpu_2_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_2_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_3_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_3_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_3_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_3_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_3_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_3_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_3_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_3_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_3_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_3_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_3_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_3_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_3_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_3_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_3_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_3_data_master_read),                                               //                          .read
		.av_readdata           (cpu_3_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_3_data_master_write),                                              //                          .write
		.av_writedata          (cpu_3_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_3_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_2_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_2_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_2_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_2_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_2_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_2_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_2_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_2_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_2_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_2_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_2_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_2_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_2_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_2_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_2_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_2_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_2_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_3_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_3_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_3_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_3_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_3_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_3_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_3_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_3_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_3_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_3_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_3_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_3_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_3_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_3_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_3_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_3_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_3_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_4_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_4_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_4_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_4_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_4_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_4_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_4_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_4_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_4_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_4_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_4_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_4_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_4_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_4_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_4_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_4_data_master_read),                                               //                          .read
		.av_readdata           (cpu_4_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_4_data_master_write),                                              //                          .write
		.av_writedata          (cpu_4_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_4_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_4_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_4_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_4_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_4_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_4_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_4_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_4_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_4_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_4_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_4_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_4_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_4_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_4_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_4_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_4_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_4_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_4_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_5_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_5_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_5_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_5_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_5_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_5_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_5_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_5_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_5_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_5_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_5_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_5_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_5_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_5_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_5_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_5_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_5_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_0_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_controller_s1_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_015_reset_out_reset),                                             //                    reset.reset
		.uav_address           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_controller_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_controller_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_controller_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_controller_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_controller_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_controller_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_controller_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_stage1_to_2_in_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                               //                    reset.reset
		.uav_address           (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_0_stage1_to_2_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_0_stage1_to_2_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_0_stage1_to_2_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                 //              (terminated)
		.av_read               (),                                                                                 //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                             //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_byteenable         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_chipselect         (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_stage1_to_2_in_csr_translator (
		.clk                   (clk_clk),                                                                              //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_0_stage1_to_2_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_stage1_to_2_in_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                               //                    reset.reset
		.uav_address           (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_1_stage1_to_2_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_1_stage1_to_2_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_1_stage1_to_2_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                 //              (terminated)
		.av_read               (),                                                                                 //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                             //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_byteenable         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_chipselect         (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_stage1_to_2_in_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                               //                    reset.reset
		.uav_address           (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_2_stage1_to_2_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_2_stage1_to_2_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_2_stage1_to_2_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                 //              (terminated)
		.av_read               (),                                                                                 //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                             //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_byteenable         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_chipselect         (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_stage1_to_2_in_csr_translator (
		.clk                   (clk_clk),                                                                              //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_2_stage1_to_2_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_stage1_to_2_in_csr_translator (
		.clk                   (clk_clk),                                                                              //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_1_stage1_to_2_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage1_to_4_in_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_008_reset_out_reset),                                             //                    reset.reset
		.uav_address           (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_stage1_to_4_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_stage1_to_4_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_stage1_to_4_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                           //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage1_to_4_in_csr_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_008_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_stage1_to_4_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage1_to_5_in_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_009_reset_out_reset),                                             //                    reset.reset
		.uav_address           (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_stage1_to_5_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_stage1_to_5_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_stage1_to_5_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                           //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage1_to_5_in_csr_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_009_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_stage1_to_5_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage1_to_6_in_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_010_reset_out_reset),                                             //                    reset.reset
		.uav_address           (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_stage1_to_6_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_stage1_to_6_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_stage1_to_6_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_readdata           (8'b10101101),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage1_to_6_in_csr_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_010_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_stage1_to_6_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pll_pll_slave_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pll_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pll_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pll_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pll_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pll_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) instruction_mem_5_s1_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                              //                    reset.reset
		.uav_address           (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (instruction_mem_5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (instruction_mem_5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (instruction_mem_5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (instruction_mem_5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (instruction_mem_5_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (instruction_mem_5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (instruction_mem_5_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_5_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_5_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_5_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage1_to_6_out_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_010_reset_out_reset),                                              //                    reset.reset
		.uav_address           (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_stage1_to_6_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_stage1_to_6_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_stage1_to_6_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                //              (terminated)
		.av_write              (),                                                                                //              (terminated)
		.av_writedata          (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage5_to_6_out_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_014_reset_out_reset),                                              //                    reset.reset
		.uav_address           (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_stage5_to_6_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_stage5_to_6_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_stage5_to_6_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                //              (terminated)
		.av_write              (),                                                                                //              (terminated)
		.av_writedata          (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage5_to_6_in_csr_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_014_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_stage5_to_6_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) instruction_mem_1_s1_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                              //                    reset.reset
		.uav_address           (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (instruction_mem_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (instruction_mem_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (instruction_mem_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (instruction_mem_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (instruction_mem_1_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (instruction_mem_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (instruction_mem_1_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_1_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_1_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_1_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_stage1_to_2_out_translator (
		.clk                   (clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                                //                    reset.reset
		.uav_address           (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_0_stage1_to_2_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_0_stage1_to_2_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_0_stage1_to_2_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                  //              (terminated)
		.av_write              (),                                                                                  //              (terminated)
		.av_writedata          (),                                                                                  //              (terminated)
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_chipselect         (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_stage1_to_2_out_translator (
		.clk                   (clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                                //                    reset.reset
		.uav_address           (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_1_stage1_to_2_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_1_stage1_to_2_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_1_stage1_to_2_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                  //              (terminated)
		.av_write              (),                                                                                  //              (terminated)
		.av_writedata          (),                                                                                  //              (terminated)
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_chipselect         (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_stage1_to_2_out_translator (
		.clk                   (clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                                //                    reset.reset
		.uav_address           (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_2_stage1_to_2_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_2_stage1_to_2_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_2_stage1_to_2_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                  //              (terminated)
		.av_write              (),                                                                                  //              (terminated)
		.av_writedata          (),                                                                                  //              (terminated)
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_chipselect         (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage2_to_3_in_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_011_reset_out_reset),                                             //                    reset.reset
		.uav_address           (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_stage2_to_3_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_stage2_to_3_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_stage2_to_3_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                           //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage2_to_3_in_csr_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_011_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_stage2_to_3_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) instruction_mem_2_s1_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                              //                    reset.reset
		.uav_address           (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (instruction_mem_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (instruction_mem_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (instruction_mem_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (instruction_mem_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (instruction_mem_2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (instruction_mem_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (instruction_mem_2_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_2_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_2_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (cpu_2_jtag_debug_module_reset_reset),                                                      //                    reset.reset
		.uav_address           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_2_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage2_to_3_out_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_011_reset_out_reset),                                              //                    reset.reset
		.uav_address           (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_stage2_to_3_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_stage2_to_3_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_stage2_to_3_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                //              (terminated)
		.av_write              (),                                                                                //              (terminated)
		.av_writedata          (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage3_to_4_in_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_012_reset_out_reset),                                             //                    reset.reset
		.uav_address           (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_stage3_to_4_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_stage3_to_4_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_stage3_to_4_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                           //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage3_to_4_in_csr_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_012_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_stage3_to_4_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) instruction_mem_3_s1_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                              //                    reset.reset
		.uav_address           (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (instruction_mem_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (instruction_mem_3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (instruction_mem_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (instruction_mem_3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (instruction_mem_3_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (instruction_mem_3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (instruction_mem_3_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_3_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_3_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_3_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage1_to_4_out_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_008_reset_out_reset),                                              //                    reset.reset
		.uav_address           (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_stage1_to_4_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_stage1_to_4_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_stage1_to_4_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                //              (terminated)
		.av_write              (),                                                                                //              (terminated)
		.av_writedata          (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage3_to_4_out_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_012_reset_out_reset),                                              //                    reset.reset
		.uav_address           (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_stage3_to_4_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_stage3_to_4_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_stage3_to_4_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                //              (terminated)
		.av_write              (),                                                                                //              (terminated)
		.av_writedata          (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage4_to_5_in_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_013_reset_out_reset),                                             //                    reset.reset
		.uav_address           (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_stage4_to_5_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_stage4_to_5_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_stage4_to_5_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                           //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage4_to_5_in_csr_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_013_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_stage4_to_5_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) instruction_mem_4_s1_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                              //                    reset.reset
		.uav_address           (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (instruction_mem_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (instruction_mem_4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (instruction_mem_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (instruction_mem_4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (instruction_mem_4_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (instruction_mem_4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (instruction_mem_4_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_4_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_4_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_4_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage1_to_5_out_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_009_reset_out_reset),                                              //                    reset.reset
		.uav_address           (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_stage1_to_5_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_stage1_to_5_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_stage1_to_5_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                //              (terminated)
		.av_write              (),                                                                                //              (terminated)
		.av_writedata          (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage4_to_5_out_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_013_reset_out_reset),                                              //                    reset.reset
		.uav_address           (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_stage4_to_5_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_stage4_to_5_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_stage4_to_5_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                //              (terminated)
		.av_write              (),                                                                                //              (terminated)
		.av_writedata          (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_stage5_to_6_in_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_014_reset_out_reset),                                             //                    reset.reset
		.uav_address           (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_stage5_to_6_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_stage5_to_6_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_stage5_to_6_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                           //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                 //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                              //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                        //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                          //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                 //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_5_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_5_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_5_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_5_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_5_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_5_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_5_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_5_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_5_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_5_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_5_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_5_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_002_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_002_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_002_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_002_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_002_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_002_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_4_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_4_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_4_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_4_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_4_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_4_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_4_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_4_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_4_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_4_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_4_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_4_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_003_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_003_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_003_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_003_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_003_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_003_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_4_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_4_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_4_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_4_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_4_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_4_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_4_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_4_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_4_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_4_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_4_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_4_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (5),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_1_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_1_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_1_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_1_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_1_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_1_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_1_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_1_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_1_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_1_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_1_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_1_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_002_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_002_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_002_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_002_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_002_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_002_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (6),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_1_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_1_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_1_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_1_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_1_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_1_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_1_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_1_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_1_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_1_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_1_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_1_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_006_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_006_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_006_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_006_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_006_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_006_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (7),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_2_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_2_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_2_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_2_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_2_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_2_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_2_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_2_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_2_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_2_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_2_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_2_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_007_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_007_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_007_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_007_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_007_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_007_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (8),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_3_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_3_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_3_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_3_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_3_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_3_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_3_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_3_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_3_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_3_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_3_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_3_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_008_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_008_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_008_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_008_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_008_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_008_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (9),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_3_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_3_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_3_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_3_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_3_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_3_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_3_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_3_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_3_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_3_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_3_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_3_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_003_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_003_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_003_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_003_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_003_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_003_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (10),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_2_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_2_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_2_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_2_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_2_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_2_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_2_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_2_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_2_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_2_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_2_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_2_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_004_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_004_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_004_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_004_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_004_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_004_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (11),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_5_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_5_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_5_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_5_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_5_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_5_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_5_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_5_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_5_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_5_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_5_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_5_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_005_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_005_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_005_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_005_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_005_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_005_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_controller_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_015_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                             //                .channel
		.rf_sink_ready           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_015_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                 //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                            //                .channel
		.rf_sink_ready           (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                                   //                .channel
		.rf_sink_ready           (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                            //                .channel
		.rf_sink_ready           (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                            //                .channel
		.rf_sink_ready           (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                                   //                .channel
		.rf_sink_ready           (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                                   //                .channel
		.rf_sink_ready           (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_008_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_008_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_008_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_011_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_011_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_011_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_011_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_011_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_011_src_channel),                                                                 //                .channel
		.rf_sink_ready           (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_008_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_009_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_009_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_009_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_013_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_013_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_013_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_013_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_013_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_013_src_channel),                                                                 //                .channel
		.rf_sink_ready           (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_009_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (56),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (36),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (37),
		.PKT_TRANS_POSTED          (38),
		.PKT_TRANS_WRITE           (39),
		.PKT_TRANS_READ            (40),
		.PKT_TRANS_LOCK            (41),
		.PKT_SRC_ID_H              (63),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (64),
		.PKT_BURSTWRAP_H           (48),
		.PKT_BURSTWRAP_L           (46),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (43),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (51),
		.PKT_BURST_SIZE_L          (49),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_010_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                              //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                              //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                               //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                        //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                            //                .channel
		.rf_sink_ready           (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_010_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_010_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_015_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_015_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_015_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_015_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_015_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_015_src_channel),                                                                 //                .channel
		.rf_sink_ready           (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_010_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                   //                .channel
		.rf_sink_ready           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) instruction_mem_5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_017_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_017_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_017_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_017_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_017_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_017_src_channel),                                                              //                .channel
		.rf_sink_ready           (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_018_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_018_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_018_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_018_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_018_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_018_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src4_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src4_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_002_src4_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src4_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src4_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src4_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src5_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src5_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src5_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src5_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src5_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src5_channel),                                                 //                .channel
		.rf_sink_ready           (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (56),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (36),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (37),
		.PKT_TRANS_POSTED          (38),
		.PKT_TRANS_WRITE           (39),
		.PKT_TRANS_READ            (40),
		.PKT_TRANS_LOCK            (41),
		.PKT_SRC_ID_H              (63),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (64),
		.PKT_BURSTWRAP_H           (48),
		.PKT_BURSTWRAP_L           (46),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (43),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (51),
		.PKT_BURST_SIZE_L          (49),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_010_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                           //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                           //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                            //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                     //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_010_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_014_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src7_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src7_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_002_src7_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src7_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src7_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src7_channel),                                                           //                .channel
		.rf_sink_ready           (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_014_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_014_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_023_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_023_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_023_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_023_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_023_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_023_src_channel),                                                                 //                .channel
		.rf_sink_ready           (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_014_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_013_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_024_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_024_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_024_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_024_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_024_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_024_src_channel),                                                                 //                .channel
		.rf_sink_ready           (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_013_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) instruction_mem_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_025_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_025_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_025_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_025_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_025_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_025_src_channel),                                                              //                .channel
		.rf_sink_ready           (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_026_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_026_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_026_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_026_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_026_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_026_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src6_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src6_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_003_src6_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src6_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src6_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src6_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src7_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src7_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_003_src7_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src7_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src7_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src7_channel),                                                 //                .channel
		.rf_sink_ready           (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_009_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src8_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src8_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_003_src8_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src8_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src8_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src8_channel),                                                           //                .channel
		.rf_sink_ready           (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_009_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_013_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src9_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src9_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_003_src9_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src9_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src9_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src9_channel),                                                           //                .channel
		.rf_sink_ready           (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_013_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_014_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src10_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src10_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_003_src10_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src10_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src10_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src10_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_014_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) instruction_mem_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_032_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_032_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_032_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_032_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_032_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_032_src_channel),                                                              //                .channel
		.rf_sink_ready           (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_033_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_033_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_033_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_033_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_033_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_033_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src6_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src6_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_006_src6_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src6_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src6_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src6_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src7_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src7_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_006_src7_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src7_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src7_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src7_channel),                                                 //                .channel
		.rf_sink_ready           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src8_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src8_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_006_src8_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src8_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src8_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src8_channel),                                                             //                .channel
		.rf_sink_ready           (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src9_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src9_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_006_src9_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src9_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src9_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src9_channel),                                                             //                .channel
		.rf_sink_ready           (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src10_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src10_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_006_src10_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src10_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src10_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src10_channel),                                                            //                .channel
		.rf_sink_ready           (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_011_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src11_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src11_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_006_src11_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src11_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src11_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src11_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_011_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_011_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_040_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_040_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_040_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_040_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_040_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_040_src_channel),                                                                 //                .channel
		.rf_sink_ready           (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_011_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) instruction_mem_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_041_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_041_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_041_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_041_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_041_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_041_src_channel),                                                              //                .channel
		.rf_sink_ready           (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_042_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_042_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_042_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_042_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_042_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_042_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (cpu_2_jtag_debug_module_reset_reset),                                                                //       clk_reset.reset
		.m0_address              (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src4_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src4_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_007_src4_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src4_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src4_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src4_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (cpu_2_jtag_debug_module_reset_reset),                                                                // clk_reset.reset
		.in_data           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src5_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src5_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_007_src5_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src5_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src5_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src5_channel),                                                 //                .channel
		.rf_sink_ready           (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_011_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src6_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src6_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_007_src6_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src6_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src6_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src6_channel),                                                           //                .channel
		.rf_sink_ready           (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_011_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_012_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src7_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src7_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_007_src7_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src7_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src7_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src7_channel),                                                          //                .channel
		.rf_sink_ready           (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_012_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_012_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_047_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_047_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_047_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_047_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_047_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_047_src_channel),                                                                 //                .channel
		.rf_sink_ready           (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_012_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) instruction_mem_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_048_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_048_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_048_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_048_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_048_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_048_src_channel),                                                              //                .channel
		.rf_sink_ready           (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_049_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_049_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_049_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_049_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_049_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_049_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src6_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src6_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_008_src6_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src6_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src6_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src6_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src7_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src7_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_008_src7_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src7_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src7_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src7_channel),                                                 //                .channel
		.rf_sink_ready           (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_008_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src8_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src8_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_008_src8_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src8_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src8_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src8_channel),                                                           //                .channel
		.rf_sink_ready           (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_008_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_012_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src9_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src9_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_008_src9_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src9_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src9_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src9_channel),                                                           //                .channel
		.rf_sink_ready           (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_012_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (55),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_013_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src10_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src10_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_008_src10_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src10_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src10_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src10_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_013_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	SoC_addr_router addr_router (
		.sink_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	SoC_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_002 addr_router_002 (
		.sink_ready         (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                     //          .valid
		.src_data           (addr_router_002_src_data),                                                      //          .data
		.src_channel        (addr_router_002_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_003 addr_router_003 (
		.sink_ready         (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                     //          .valid
		.src_data           (addr_router_003_src_data),                                                      //          .data
		.src_channel        (addr_router_003_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_004 addr_router_004 (
		.sink_ready         (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                            //          .valid
		.src_data           (addr_router_004_src_data),                                                             //          .data
		.src_channel        (addr_router_004_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_addr_router_005 addr_router_005 (
		.sink_ready         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                            //          .valid
		.src_data           (addr_router_005_src_data),                                                             //          .data
		.src_channel        (addr_router_005_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_addr_router_006 addr_router_006 (
		.sink_ready         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                     //          .valid
		.src_data           (addr_router_006_src_data),                                                      //          .data
		.src_channel        (addr_router_006_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_007 addr_router_007 (
		.sink_ready         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_007_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_007_src_valid),                                                     //          .valid
		.src_data           (addr_router_007_src_data),                                                      //          .data
		.src_channel        (addr_router_007_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_007_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_007_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_008 addr_router_008 (
		.sink_ready         (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_008_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_008_src_valid),                                                     //          .valid
		.src_data           (addr_router_008_src_data),                                                      //          .data
		.src_channel        (addr_router_008_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_008_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_008_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_009 addr_router_009 (
		.sink_ready         (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_009_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_009_src_valid),                                                            //          .valid
		.src_data           (addr_router_009_src_data),                                                             //          .data
		.src_channel        (addr_router_009_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_009_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_009_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_addr_router_010 addr_router_010 (
		.sink_ready         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_010_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_010_src_valid),                                                            //          .valid
		.src_data           (addr_router_010_src_data),                                                             //          .data
		.src_channel        (addr_router_010_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_010_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_010_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_addr_router_011 addr_router_011 (
		.sink_ready         (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_011_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_011_src_valid),                                                            //          .valid
		.src_data           (addr_router_011_src_data),                                                             //          .data
		.src_channel        (addr_router_011_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_011_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_011_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router id_router (
		.sink_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	SoC_id_router_001 id_router_001 (
		.sink_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_015_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                        //       src.ready
		.src_valid          (id_router_001_src_valid),                                                        //          .valid
		.src_data           (id_router_001_src_data),                                                         //          .data
		.src_channel        (id_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	SoC_id_router_002 id_router_002 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                               //       src.ready
		.src_valid          (id_router_002_src_valid),                                               //          .valid
		.src_data           (id_router_002_src_data),                                                //          .data
		.src_channel        (id_router_002_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_002 id_router_003 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                  //          .valid
		.src_data           (id_router_003_src_data),                                                                   //          .data
		.src_channel        (id_router_003_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_002 id_router_004 (
		.sink_ready         (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                          //       src.ready
		.src_valid          (id_router_004_src_valid),                                                          //          .valid
		.src_data           (id_router_004_src_data),                                                           //          .data
		.src_channel        (id_router_004_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                     //          .endofpacket
	);

	SoC_id_router_005 id_router_005 (
		.sink_ready         (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                              //       src.ready
		.src_valid          (id_router_005_src_valid),                                                              //          .valid
		.src_data           (id_router_005_src_data),                                                               //          .data
		.src_channel        (id_router_005_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                         //          .endofpacket
	);

	SoC_id_router_002 id_router_006 (
		.sink_ready         (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                          //       src.ready
		.src_valid          (id_router_006_src_valid),                                                          //          .valid
		.src_data           (id_router_006_src_data),                                                           //          .data
		.src_channel        (id_router_006_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                     //          .endofpacket
	);

	SoC_id_router_002 id_router_007 (
		.sink_ready         (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_stage1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                          //       src.ready
		.src_valid          (id_router_007_src_valid),                                                          //          .valid
		.src_data           (id_router_007_src_data),                                                           //          .data
		.src_channel        (id_router_007_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                     //          .endofpacket
	);

	SoC_id_router_005 id_router_008 (
		.sink_ready         (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                              //       src.ready
		.src_valid          (id_router_008_src_valid),                                                              //          .valid
		.src_data           (id_router_008_src_data),                                                               //          .data
		.src_channel        (id_router_008_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                         //          .endofpacket
	);

	SoC_id_router_005 id_router_009 (
		.sink_ready         (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_stage1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                              //       src.ready
		.src_valid          (id_router_009_src_valid),                                                              //          .valid
		.src_data           (id_router_009_src_data),                                                               //          .data
		.src_channel        (id_router_009_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                         //          .endofpacket
	);

	SoC_id_router_002 id_router_010 (
		.sink_ready         (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage1_to_4_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                        //       src.ready
		.src_valid          (id_router_010_src_valid),                                                        //          .valid
		.src_data           (id_router_010_src_data),                                                         //          .data
		.src_channel        (id_router_010_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                   //          .endofpacket
	);

	SoC_id_router_011 id_router_011 (
		.sink_ready         (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage1_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                            //       src.ready
		.src_valid          (id_router_011_src_valid),                                                            //          .valid
		.src_data           (id_router_011_src_data),                                                             //          .data
		.src_channel        (id_router_011_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_002 id_router_012 (
		.sink_ready         (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage1_to_5_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                        //       src.ready
		.src_valid          (id_router_012_src_valid),                                                        //          .valid
		.src_data           (id_router_012_src_data),                                                         //          .data
		.src_channel        (id_router_012_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                   //          .endofpacket
	);

	SoC_id_router_013 id_router_013 (
		.sink_ready         (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage1_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                            //       src.ready
		.src_valid          (id_router_013_src_valid),                                                            //          .valid
		.src_data           (id_router_013_src_data),                                                             //          .data
		.src_channel        (id_router_013_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_014 id_router_014 (
		.sink_ready         (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage1_to_6_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                        //       src.ready
		.src_valid          (id_router_014_src_valid),                                                        //          .valid
		.src_data           (id_router_014_src_data),                                                         //          .data
		.src_channel        (id_router_014_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                   //          .endofpacket
	);

	SoC_id_router_015 id_router_015 (
		.sink_ready         (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage1_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                            //       src.ready
		.src_valid          (id_router_015_src_valid),                                                            //          .valid
		.src_data           (id_router_015_src_data),                                                             //          .data
		.src_channel        (id_router_015_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_002 id_router_016 (
		.sink_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                  //       src.ready
		.src_valid          (id_router_016_src_valid),                                                  //          .valid
		.src_data           (id_router_016_src_data),                                                   //          .data
		.src_channel        (id_router_016_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_017 id_router_017 (
		.sink_ready         (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (instruction_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                         //       src.ready
		.src_valid          (id_router_017_src_valid),                                                         //          .valid
		.src_data           (id_router_017_src_data),                                                          //          .data
		.src_channel        (id_router_017_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_017 id_router_018 (
		.sink_ready         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                            //       src.ready
		.src_valid          (id_router_018_src_valid),                                                            //          .valid
		.src_data           (id_router_018_src_data),                                                             //          .data
		.src_channel        (id_router_018_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_019 id_router_019 (
		.sink_ready         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_019_src_valid),                                                                  //          .valid
		.src_data           (id_router_019_src_data),                                                                   //          .data
		.src_channel        (id_router_019_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_019 id_router_020 (
		.sink_ready         (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                               //       src.ready
		.src_valid          (id_router_020_src_valid),                                               //          .valid
		.src_data           (id_router_020_src_data),                                                //          .data
		.src_channel        (id_router_020_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_021 id_router_021 (
		.sink_ready         (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage1_to_6_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                         //       src.ready
		.src_valid          (id_router_021_src_valid),                                                         //          .valid
		.src_data           (id_router_021_src_data),                                                          //          .data
		.src_channel        (id_router_021_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_019 id_router_022 (
		.sink_ready         (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage5_to_6_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                         //       src.ready
		.src_valid          (id_router_022_src_valid),                                                         //          .valid
		.src_data           (id_router_022_src_data),                                                          //          .data
		.src_channel        (id_router_022_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_023 id_router_023 (
		.sink_ready         (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage5_to_6_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                                            //       src.ready
		.src_valid          (id_router_023_src_valid),                                                            //          .valid
		.src_data           (id_router_023_src_data),                                                             //          .data
		.src_channel        (id_router_023_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_024 id_router_024 (
		.sink_ready         (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage4_to_5_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                                            //       src.ready
		.src_valid          (id_router_024_src_valid),                                                            //          .valid
		.src_data           (id_router_024_src_data),                                                             //          .data
		.src_channel        (id_router_024_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_025 id_router_025 (
		.sink_ready         (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (instruction_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                         //       src.ready
		.src_valid          (id_router_025_src_valid),                                                         //          .valid
		.src_data           (id_router_025_src_data),                                                          //          .data
		.src_channel        (id_router_025_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_025 id_router_026 (
		.sink_ready         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                            //       src.ready
		.src_valid          (id_router_026_src_valid),                                                            //          .valid
		.src_data           (id_router_026_src_data),                                                             //          .data
		.src_channel        (id_router_026_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_027 id_router_027 (
		.sink_ready         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_027_src_valid),                                                                  //          .valid
		.src_data           (id_router_027_src_data),                                                                   //          .data
		.src_channel        (id_router_027_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_027 id_router_028 (
		.sink_ready         (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                               //       src.ready
		.src_valid          (id_router_028_src_valid),                                               //          .valid
		.src_data           (id_router_028_src_data),                                                //          .data
		.src_channel        (id_router_028_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_027 id_router_029 (
		.sink_ready         (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage1_to_5_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                                         //       src.ready
		.src_valid          (id_router_029_src_valid),                                                         //          .valid
		.src_data           (id_router_029_src_data),                                                          //          .data
		.src_channel        (id_router_029_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_027 id_router_030 (
		.sink_ready         (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage4_to_5_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                                         //       src.ready
		.src_valid          (id_router_030_src_valid),                                                         //          .valid
		.src_data           (id_router_030_src_data),                                                          //          .data
		.src_channel        (id_router_030_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_027 id_router_031 (
		.sink_ready         (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage5_to_6_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_031_src_ready),                                                        //       src.ready
		.src_valid          (id_router_031_src_valid),                                                        //          .valid
		.src_data           (id_router_031_src_data),                                                         //          .data
		.src_channel        (id_router_031_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_031_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_031_src_endofpacket)                                                   //          .endofpacket
	);

	SoC_id_router_032 id_router_032 (
		.sink_ready         (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (instruction_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_032_src_ready),                                                         //       src.ready
		.src_valid          (id_router_032_src_valid),                                                         //          .valid
		.src_data           (id_router_032_src_data),                                                          //          .data
		.src_channel        (id_router_032_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_032_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_032_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_032 id_router_033 (
		.sink_ready         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_033_src_ready),                                                            //       src.ready
		.src_valid          (id_router_033_src_valid),                                                            //          .valid
		.src_data           (id_router_033_src_data),                                                             //          .data
		.src_channel        (id_router_033_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_033_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_033_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_034 id_router_034 (
		.sink_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_034_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_034_src_valid),                                                                  //          .valid
		.src_data           (id_router_034_src_data),                                                                   //          .data
		.src_channel        (id_router_034_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_034_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_034_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_034 id_router_035 (
		.sink_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_035_src_ready),                                               //       src.ready
		.src_valid          (id_router_035_src_valid),                                               //          .valid
		.src_data           (id_router_035_src_data),                                                //          .data
		.src_channel        (id_router_035_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_035_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_035_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_034 id_router_036 (
		.sink_ready         (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_036_src_ready),                                                           //       src.ready
		.src_valid          (id_router_036_src_valid),                                                           //          .valid
		.src_data           (id_router_036_src_data),                                                            //          .data
		.src_channel        (id_router_036_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_036_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_036_src_endofpacket)                                                      //          .endofpacket
	);

	SoC_id_router_034 id_router_037 (
		.sink_ready         (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_037_src_ready),                                                           //       src.ready
		.src_valid          (id_router_037_src_valid),                                                           //          .valid
		.src_data           (id_router_037_src_data),                                                            //          .data
		.src_channel        (id_router_037_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_037_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_037_src_endofpacket)                                                      //          .endofpacket
	);

	SoC_id_router_034 id_router_038 (
		.sink_ready         (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_stage1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_038_src_ready),                                                           //       src.ready
		.src_valid          (id_router_038_src_valid),                                                           //          .valid
		.src_data           (id_router_038_src_data),                                                            //          .data
		.src_channel        (id_router_038_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_038_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_038_src_endofpacket)                                                      //          .endofpacket
	);

	SoC_id_router_034 id_router_039 (
		.sink_ready         (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage2_to_3_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_039_src_ready),                                                        //       src.ready
		.src_valid          (id_router_039_src_valid),                                                        //          .valid
		.src_data           (id_router_039_src_data),                                                         //          .data
		.src_channel        (id_router_039_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_039_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_039_src_endofpacket)                                                   //          .endofpacket
	);

	SoC_id_router_040 id_router_040 (
		.sink_ready         (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage2_to_3_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_040_src_ready),                                                            //       src.ready
		.src_valid          (id_router_040_src_valid),                                                            //          .valid
		.src_data           (id_router_040_src_data),                                                             //          .data
		.src_channel        (id_router_040_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_040_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_040_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_041 id_router_041 (
		.sink_ready         (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (instruction_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_041_src_ready),                                                         //       src.ready
		.src_valid          (id_router_041_src_valid),                                                         //          .valid
		.src_data           (id_router_041_src_data),                                                          //          .data
		.src_channel        (id_router_041_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_041_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_041_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_041 id_router_042 (
		.sink_ready         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_042_src_ready),                                                            //       src.ready
		.src_valid          (id_router_042_src_valid),                                                            //          .valid
		.src_data           (id_router_042_src_data),                                                             //          .data
		.src_channel        (id_router_042_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_042_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_042_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_043 id_router_043 (
		.sink_ready         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (cpu_2_jtag_debug_module_reset_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_043_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_043_src_valid),                                                                  //          .valid
		.src_data           (id_router_043_src_data),                                                                   //          .data
		.src_channel        (id_router_043_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_043_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_043_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_043 id_router_044 (
		.sink_ready         (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_044_src_ready),                                               //       src.ready
		.src_valid          (id_router_044_src_valid),                                               //          .valid
		.src_data           (id_router_044_src_data),                                                //          .data
		.src_channel        (id_router_044_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_044_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_044_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_043 id_router_045 (
		.sink_ready         (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage2_to_3_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_045_src_ready),                                                         //       src.ready
		.src_valid          (id_router_045_src_valid),                                                         //          .valid
		.src_data           (id_router_045_src_data),                                                          //          .data
		.src_channel        (id_router_045_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_045_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_045_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_043 id_router_046 (
		.sink_ready         (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage3_to_4_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_046_src_ready),                                                        //       src.ready
		.src_valid          (id_router_046_src_valid),                                                        //          .valid
		.src_data           (id_router_046_src_data),                                                         //          .data
		.src_channel        (id_router_046_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_046_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_046_src_endofpacket)                                                   //          .endofpacket
	);

	SoC_id_router_047 id_router_047 (
		.sink_ready         (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage3_to_4_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_047_src_ready),                                                            //       src.ready
		.src_valid          (id_router_047_src_valid),                                                            //          .valid
		.src_data           (id_router_047_src_data),                                                             //          .data
		.src_channel        (id_router_047_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_047_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_047_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_048 id_router_048 (
		.sink_ready         (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (instruction_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_048_src_ready),                                                         //       src.ready
		.src_valid          (id_router_048_src_valid),                                                         //          .valid
		.src_data           (id_router_048_src_data),                                                          //          .data
		.src_channel        (id_router_048_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_048_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_048_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_048 id_router_049 (
		.sink_ready         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_049_src_ready),                                                            //       src.ready
		.src_valid          (id_router_049_src_valid),                                                            //          .valid
		.src_data           (id_router_049_src_data),                                                             //          .data
		.src_channel        (id_router_049_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_049_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_049_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_050 id_router_050 (
		.sink_ready         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_050_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_050_src_valid),                                                                  //          .valid
		.src_data           (id_router_050_src_data),                                                                   //          .data
		.src_channel        (id_router_050_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_050_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_050_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_050 id_router_051 (
		.sink_ready         (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_051_src_ready),                                               //       src.ready
		.src_valid          (id_router_051_src_valid),                                               //          .valid
		.src_data           (id_router_051_src_data),                                                //          .data
		.src_channel        (id_router_051_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_051_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_051_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_050 id_router_052 (
		.sink_ready         (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage1_to_4_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_052_src_ready),                                                         //       src.ready
		.src_valid          (id_router_052_src_valid),                                                         //          .valid
		.src_data           (id_router_052_src_data),                                                          //          .data
		.src_channel        (id_router_052_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_052_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_052_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_050 id_router_053 (
		.sink_ready         (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage3_to_4_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_053_src_ready),                                                         //       src.ready
		.src_valid          (id_router_053_src_valid),                                                         //          .valid
		.src_data           (id_router_053_src_data),                                                          //          .data
		.src_channel        (id_router_053_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_053_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_053_src_endofpacket)                                                    //          .endofpacket
	);

	SoC_id_router_050 id_router_054 (
		.sink_ready         (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_stage4_to_5_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_054_src_ready),                                                        //       src.ready
		.src_valid          (id_router_054_src_valid),                                                        //          .valid
		.src_data           (id_router_054_src_data),                                                         //          .data
		.src_channel        (id_router_054_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_054_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_054_src_endofpacket)                                                   //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.VALID_WIDTH               (55),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.VALID_WIDTH               (55),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_004_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_004_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_004_src_data),           //          .data
		.cmd_sink_channel       (addr_router_004_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_004_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_004_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_004_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_004_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_004_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_004_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_004_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_004_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.VALID_WIDTH               (55),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_005_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_005_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_005_src_data),           //          .data
		.cmd_sink_channel       (addr_router_005_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_005_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_005_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_005_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_005_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_005_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_005_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_005_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_005_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.VALID_WIDTH               (55),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_003 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_009_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_009_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_009_src_data),           //          .data
		.cmd_sink_channel       (addr_router_009_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_009_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_009_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_003_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_003_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_003_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_003_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_003_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_009_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_009_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_009_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_009_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_009_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_009_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_003_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_003_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_003_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_003_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_003_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_003_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_003_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.VALID_WIDTH               (55),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_004 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_010_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_010_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_010_src_data),           //          .data
		.cmd_sink_channel       (addr_router_010_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_010_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_010_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_004_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_004_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_004_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_004_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_004_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_010_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_010_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_010_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_010_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_010_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_010_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_004_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_004_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_004_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_004_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_004_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_004_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_004_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (91),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (55),
		.VALID_WIDTH               (55),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_005 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_011_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_011_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_011_src_data),           //          .data
		.cmd_sink_channel       (addr_router_011_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_011_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_011_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_005_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_005_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_005_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_005_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_005_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_011_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_011_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_011_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_011_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_011_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_011_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_005_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_005_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_005_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_005_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_005_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_005_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_005_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (36),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (56),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (43),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (51),
		.PKT_BURST_SIZE_L          (49),
		.PKT_BURST_TYPE_H          (53),
		.PKT_BURST_TYPE_L          (52),
		.PKT_BURSTWRAP_H           (48),
		.PKT_BURSTWRAP_L           (46),
		.PKT_TRANS_COMPRESSED_READ (37),
		.PKT_TRANS_WRITE           (39),
		.PKT_TRANS_READ            (40),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (55),
		.OUT_BYTE_CNT_H            (43),
		.OUT_BURSTWRAP_H           (48),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter (
		.clk                   (clk_clk),                             //       cr0.clk
		.reset                 (rst_controller_010_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (36),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (56),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (43),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (51),
		.PKT_BURST_SIZE_L          (49),
		.PKT_BURST_TYPE_H          (53),
		.PKT_BURST_TYPE_L          (52),
		.PKT_BURSTWRAP_H           (48),
		.PKT_BURSTWRAP_L           (46),
		.PKT_TRANS_COMPRESSED_READ (37),
		.PKT_TRANS_WRITE           (39),
		.PKT_TRANS_READ            (40),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (55),
		.OUT_BYTE_CNT_H            (43),
		.OUT_BURSTWRAP_H           (48),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_010_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_1_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_004 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_3_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_005 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_4_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_006 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_5_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_006_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_007 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_1_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_007_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_008 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_3_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_008_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_009 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_4_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_009_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_010 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_5_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_010_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_011 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_1_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_2_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_011_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_012 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_2_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_3_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_012_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_013 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_3_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_4_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_013_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_014 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_4_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_5_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_014_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (7),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_015 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_1_jtag_debug_module_reset_reset), // reset_in2.reset
		.reset_in3  (cpu_2_jtag_debug_module_reset_reset), // reset_in3.reset
		.reset_in4  (cpu_3_jtag_debug_module_reset_reset), // reset_in4.reset
		.reset_in5  (cpu_4_jtag_debug_module_reset_reset), // reset_in5.reset
		.reset_in6  (cpu_5_jtag_debug_module_reset_reset), // reset_in6.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_015_reset_out_reset),  // reset_out.reset
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	SoC_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_002_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_002_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_002_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_002_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_002_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_002_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_002_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_002_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_002_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_002_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_002_src5_endofpacket),   //          .endofpacket
		.src6_ready         (cmd_xbar_demux_002_src6_ready),         //      src6.ready
		.src6_valid         (cmd_xbar_demux_002_src6_valid),         //          .valid
		.src6_data          (cmd_xbar_demux_002_src6_data),          //          .data
		.src6_channel       (cmd_xbar_demux_002_src6_channel),       //          .channel
		.src6_startofpacket (cmd_xbar_demux_002_src6_startofpacket), //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_002_src6_endofpacket),   //          .endofpacket
		.src7_ready         (cmd_xbar_demux_002_src7_ready),         //      src7.ready
		.src7_valid         (cmd_xbar_demux_002_src7_valid),         //          .valid
		.src7_data          (cmd_xbar_demux_002_src7_data),          //          .data
		.src7_channel       (cmd_xbar_demux_002_src7_channel),       //          .channel
		.src7_startofpacket (cmd_xbar_demux_002_src7_startofpacket), //          .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_002_src7_endofpacket),   //          .endofpacket
		.src8_ready         (cmd_xbar_demux_002_src8_ready),         //      src8.ready
		.src8_valid         (cmd_xbar_demux_002_src8_valid),         //          .valid
		.src8_data          (cmd_xbar_demux_002_src8_data),          //          .data
		.src8_channel       (cmd_xbar_demux_002_src8_channel),       //          .channel
		.src8_startofpacket (cmd_xbar_demux_002_src8_startofpacket), //          .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_002_src8_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_003_src_ready),              //      sink.ready
		.sink_channel        (addr_router_003_src_channel),            //          .channel
		.sink_data           (addr_router_003_src_data),               //          .data
		.sink_startofpacket  (addr_router_003_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_003_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_003_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_003_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_003_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_003_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_003_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_003_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_003_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_003_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_003_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_003_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_003_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_003_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_003_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_003_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_003_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_003_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_003_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_003_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_003_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_003_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_003_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_003_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_003_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_003_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_003_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_003_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_003_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_003_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_003_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_003_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_003_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_003_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_003_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_003_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_003_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_003_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_003_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_003_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_003_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_003_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_003_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_003_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_003_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_003_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_003_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_003_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_003_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_003_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_003_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_003_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_003_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_003_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_003_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_003_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_003_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_003_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_003_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_003_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_003_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_003_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_003_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_003_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_003_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_003_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_003_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_003_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_003_src10_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_004_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_004_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_004_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_004_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_004_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_004_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_004_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_004_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_004_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_004_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_004_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_004_src2_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_004 cmd_xbar_demux_005 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_005_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_005_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_005_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_005_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_005_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_005_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_005_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_005_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_005_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_005_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_005_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_005_src2_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_006 cmd_xbar_demux_006 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_006_src_ready),              //      sink.ready
		.sink_channel        (addr_router_006_src_channel),            //          .channel
		.sink_data           (addr_router_006_src_data),               //          .data
		.sink_startofpacket  (addr_router_006_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_006_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_006_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_006_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_006_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_006_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_006_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_006_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_006_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_006_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_006_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_006_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_006_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_006_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_006_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_006_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_006_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_006_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_006_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_006_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_006_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_006_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_006_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_006_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_006_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_006_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_006_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_006_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_006_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_006_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_006_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_006_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_006_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_006_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_006_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_006_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_006_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_006_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_006_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_006_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_006_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_006_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_006_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_006_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_006_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_006_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_006_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_006_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_006_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_006_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_006_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_006_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_006_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_006_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_006_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_006_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_006_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_006_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_006_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_006_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_006_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_006_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_006_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_006_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_006_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_006_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_006_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_006_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_006_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_006_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_006_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_006_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_006_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_006_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_006_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_006_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_006_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_006_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_006_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_006_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_006_src12_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_002 cmd_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_007_src_ready),             //      sink.ready
		.sink_channel       (addr_router_007_src_channel),           //          .channel
		.sink_data          (addr_router_007_src_data),              //          .data
		.sink_startofpacket (addr_router_007_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_007_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_007_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_007_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_007_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_007_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_007_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_007_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_007_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_007_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_007_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_007_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_007_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_007_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_007_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_007_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_007_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_007_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_007_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_007_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_007_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_007_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_007_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_007_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_007_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_007_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_007_src5_endofpacket),   //          .endofpacket
		.src6_ready         (cmd_xbar_demux_007_src6_ready),         //      src6.ready
		.src6_valid         (cmd_xbar_demux_007_src6_valid),         //          .valid
		.src6_data          (cmd_xbar_demux_007_src6_data),          //          .data
		.src6_channel       (cmd_xbar_demux_007_src6_channel),       //          .channel
		.src6_startofpacket (cmd_xbar_demux_007_src6_startofpacket), //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_007_src6_endofpacket),   //          .endofpacket
		.src7_ready         (cmd_xbar_demux_007_src7_ready),         //      src7.ready
		.src7_valid         (cmd_xbar_demux_007_src7_valid),         //          .valid
		.src7_data          (cmd_xbar_demux_007_src7_data),          //          .data
		.src7_channel       (cmd_xbar_demux_007_src7_channel),       //          .channel
		.src7_startofpacket (cmd_xbar_demux_007_src7_startofpacket), //          .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_007_src7_endofpacket),   //          .endofpacket
		.src8_ready         (cmd_xbar_demux_007_src8_ready),         //      src8.ready
		.src8_valid         (cmd_xbar_demux_007_src8_valid),         //          .valid
		.src8_data          (cmd_xbar_demux_007_src8_data),          //          .data
		.src8_channel       (cmd_xbar_demux_007_src8_channel),       //          .channel
		.src8_startofpacket (cmd_xbar_demux_007_src8_startofpacket), //          .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_007_src8_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_003 cmd_xbar_demux_008 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_008_src_ready),              //      sink.ready
		.sink_channel        (addr_router_008_src_channel),            //          .channel
		.sink_data           (addr_router_008_src_data),               //          .data
		.sink_startofpacket  (addr_router_008_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_008_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_008_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_008_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_008_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_008_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_008_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_008_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_008_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_008_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_008_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_008_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_008_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_008_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_008_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_008_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_008_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_008_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_008_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_008_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_008_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_008_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_008_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_008_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_008_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_008_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_008_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_008_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_008_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_008_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_008_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_008_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_008_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_008_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_008_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_008_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_008_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_008_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_008_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_008_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_008_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_008_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_008_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_008_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_008_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_008_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_008_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_008_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_008_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_008_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_008_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_008_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_008_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_008_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_008_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_008_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_008_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_008_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_008_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_008_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_008_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_008_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_008_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_008_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_008_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_008_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_008_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_008_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_008_src10_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_004 cmd_xbar_demux_009 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_003_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_003_cmd_src_channel),           //           .channel
		.sink_data          (limiter_003_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_003_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_003_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_003_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_009_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_009_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_009_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_009_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_009_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_009_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_009_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_009_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_009_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_009_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_009_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_009_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_009_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_009_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_009_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_009_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_009_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_009_src2_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_004 cmd_xbar_demux_010 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_004_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_004_cmd_src_channel),           //           .channel
		.sink_data          (limiter_004_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_004_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_004_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_004_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_010_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_010_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_010_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_010_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_010_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_010_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_010_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_010_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_010_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_010_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_010_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_010_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_010_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_010_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_010_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_010_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_010_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_010_src2_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_004 cmd_xbar_demux_011 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_005_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_005_cmd_src_channel),           //           .channel
		.sink_data          (limiter_005_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_005_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_005_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_005_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_011_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_011_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_011_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_011_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_011_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_011_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_011_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_011_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_011_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_011_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_011_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_011_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_011_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_011_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_011_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_011_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_011_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_011_src2_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_015_reset_out_reset),    // clk_reset.reset
		.src_ready            (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data             (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel          (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (cmd_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (cmd_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (cmd_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (cmd_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (cmd_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (cmd_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (cmd_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (cmd_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (cmd_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (cmd_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (cmd_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (cmd_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (cmd_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (cmd_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (cmd_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (cmd_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (cmd_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (cmd_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (cmd_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (cmd_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (cmd_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (cmd_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (cmd_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (cmd_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (cmd_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (cmd_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (cmd_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (cmd_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (cmd_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (cmd_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (cmd_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (cmd_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (cmd_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (cmd_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (cmd_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (cmd_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (cmd_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (cmd_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (cmd_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (cmd_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (cmd_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (cmd_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (cmd_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (cmd_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (cmd_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src5_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_006_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_006_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_006_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_006_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_008 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src8_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src8_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_006_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_006_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_006_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_006_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_006_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_006_src2_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_009 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src9_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src9_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src9_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src9_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src9_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_006_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_006_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_006_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_006_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_006_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_006_src3_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_011 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_008_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_011_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_011_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_011_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_011_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_011_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_011_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src11_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_008_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_008_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_008_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_008_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_008_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_008_src1_endofpacket)     //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_013 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_009_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_013_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_013_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_013_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_013_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_013_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_013_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src13_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_003_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)     //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_015 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_010_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_015_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_015_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_015_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_015_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_015_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_015_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src15_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket)     //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_017 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_017_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_017_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_017_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_017_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_017_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_017_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src2_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_011_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_011_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_011_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_011_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_011_src1_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_018 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_018_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_018_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_018_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_018_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_018_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_018_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src3_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_011_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_011_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_011_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_011_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_011_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_011_src2_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_023 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_014_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_023_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_023_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_023_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_023_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_023_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_023_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src8_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src8_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src8_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src8_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src8_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src8_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src2_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_024 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_013_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_024_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_024_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_024_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_024_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_024_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_024_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src3_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src3_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src3_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src3_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_008_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_008_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_008_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_008_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_008_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_008_src2_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_025 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_025_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_025_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_025_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_025_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_025_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_025_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src4_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src4_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src4_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src4_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src4_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src4_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_004_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_004_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_004_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_004_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_026 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_026_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_026_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_026_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_026_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_026_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_026_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src5_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src5_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src5_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src5_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src5_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src5_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_004_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_004_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_004_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_004_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_004_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_004_src2_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_032 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_032_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_032_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_032_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_032_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_032_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_032_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_005_src1_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_005_src1_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_005_src1_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_005_src1_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_006_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_006_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_006_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_006_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_006_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_006_src4_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_033 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_033_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_033_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_033_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_033_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_033_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_033_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_005_src2_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_005_src2_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_005_src2_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_005_src2_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_005_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_005_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_006_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_006_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_006_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_006_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_006_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_006_src5_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_040 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_011_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_040_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_040_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_040_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_040_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_040_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_040_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_006_src12_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_006_src12_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_006_src12_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_006_src12_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_006_src12_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_006_src12_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_007_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_007_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_007_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_007_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_007_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_007_src1_endofpacket)     //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_041 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_041_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_041_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_041_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_041_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_041_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_041_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_007_src2_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_007_src2_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_007_src2_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_007_src2_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_007_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_007_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_010_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_010_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_010_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_010_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_010_src1_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_042 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_042_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_042_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_042_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_042_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_042_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_042_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_007_src3_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_007_src3_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_007_src3_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_007_src3_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_007_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_007_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_010_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_010_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_010_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_010_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_010_src2_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_047 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_012_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_047_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_047_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_047_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_047_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_047_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_047_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_007_src8_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_007_src8_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_007_src8_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_007_src8_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_007_src8_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_007_src8_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_008_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_008_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_008_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_008_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_008_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_008_src3_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_048 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_048_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_048_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_048_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_048_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_048_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_048_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_008_src4_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_008_src4_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_008_src4_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_008_src4_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_008_src4_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_008_src4_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_049 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_049_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_049_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_049_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_049_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_049_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_049_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_008_src5_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_008_src5_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_008_src5_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_008_src5_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_008_src5_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_008_src5_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src2_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_015_reset_out_reset),     // clk_reset.reset
		.sink_ready          (id_router_001_src_ready),                //      sink.ready
		.sink_channel        (id_router_001_src_channel),              //          .channel
		.sink_data           (id_router_001_src_data),                 //          .data
		.sink_startofpacket  (id_router_001_src_startofpacket),        //          .startofpacket
		.sink_endofpacket    (id_router_001_src_endofpacket),          //          .endofpacket
		.sink_valid          (id_router_001_src_valid),                //          .valid
		.src0_ready          (rsp_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (rsp_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (rsp_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (rsp_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (rsp_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (rsp_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (rsp_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (rsp_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (rsp_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (rsp_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (rsp_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (rsp_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (rsp_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (rsp_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (rsp_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (rsp_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (rsp_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (rsp_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (rsp_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (rsp_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (rsp_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (rsp_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (rsp_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (rsp_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (rsp_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (rsp_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (rsp_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (rsp_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (rsp_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (rsp_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (rsp_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (rsp_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (rsp_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (rsp_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (rsp_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (rsp_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (rsp_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (rsp_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (rsp_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (rsp_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (rsp_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (rsp_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (rsp_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (rsp_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (rsp_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (rsp_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (rsp_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (rsp_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (rsp_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (rsp_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (rsp_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (rsp_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (rsp_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (rsp_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (rsp_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (rsp_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (rsp_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (rsp_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (rsp_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (rsp_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (rsp_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (rsp_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (rsp_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (rsp_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (rsp_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (rsp_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (rsp_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (rsp_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (rsp_xbar_demux_001_src11_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_011_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_011_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_011_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_011_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_011_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_013_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_013_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_014 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_015 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_015_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_015_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_016 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_017 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_017_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_017_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_017_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_017_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_017_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_017_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_018 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_018_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_018_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_018_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_018_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_018_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_018_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_019 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_020 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_021 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_022 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_023 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_023_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_023_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_023_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_023_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_023_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_023_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_024 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_024_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_024_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_024_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_024_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_024_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_024_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_025 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_025_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_025_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_025_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_025_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_025_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_025_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_026 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_026_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_026_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_026_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_026_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_026_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_026_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_027 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_028 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_029 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_029_src_ready),               //      sink.ready
		.sink_channel       (id_router_029_src_channel),             //          .channel
		.sink_data          (id_router_029_src_data),                //          .data
		.sink_startofpacket (id_router_029_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_029_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_029_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_030 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_030_src_ready),               //      sink.ready
		.sink_channel       (id_router_030_src_channel),             //          .channel
		.sink_data          (id_router_030_src_data),                //          .data
		.sink_startofpacket (id_router_030_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_030_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_030_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_031 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_031_src_ready),               //      sink.ready
		.sink_channel       (id_router_031_src_channel),             //          .channel
		.sink_data          (id_router_031_src_data),                //          .data
		.sink_startofpacket (id_router_031_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_031_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_031_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_031_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_032 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_032_src_ready),               //      sink.ready
		.sink_channel       (id_router_032_src_channel),             //          .channel
		.sink_data          (id_router_032_src_data),                //          .data
		.sink_startofpacket (id_router_032_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_032_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_032_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_032_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_032_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_032_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_032_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_032_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_032_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_032_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_032_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_033 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_033_src_ready),               //      sink.ready
		.sink_channel       (id_router_033_src_channel),             //          .channel
		.sink_data          (id_router_033_src_data),                //          .data
		.sink_startofpacket (id_router_033_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_033_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_033_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_033_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_033_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_033_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_033_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_033_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_033_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_033_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_033_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_034 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_034_src_ready),               //      sink.ready
		.sink_channel       (id_router_034_src_channel),             //          .channel
		.sink_data          (id_router_034_src_data),                //          .data
		.sink_startofpacket (id_router_034_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_034_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_034_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_034_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_034_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_035 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_035_src_ready),               //      sink.ready
		.sink_channel       (id_router_035_src_channel),             //          .channel
		.sink_data          (id_router_035_src_data),                //          .data
		.sink_startofpacket (id_router_035_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_035_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_035_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_035_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_035_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_036 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_036_src_ready),               //      sink.ready
		.sink_channel       (id_router_036_src_channel),             //          .channel
		.sink_data          (id_router_036_src_data),                //          .data
		.sink_startofpacket (id_router_036_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_036_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_036_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_036_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_037 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_037_src_ready),               //      sink.ready
		.sink_channel       (id_router_037_src_channel),             //          .channel
		.sink_data          (id_router_037_src_data),                //          .data
		.sink_startofpacket (id_router_037_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_037_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_037_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_037_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_037_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_038 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_038_src_ready),               //      sink.ready
		.sink_channel       (id_router_038_src_channel),             //          .channel
		.sink_data          (id_router_038_src_data),                //          .data
		.sink_startofpacket (id_router_038_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_038_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_038_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_038_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_038_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_038_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_038_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_038_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_039 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_039_src_ready),               //      sink.ready
		.sink_channel       (id_router_039_src_channel),             //          .channel
		.sink_data          (id_router_039_src_data),                //          .data
		.sink_startofpacket (id_router_039_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_039_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_039_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_039_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_039_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_039_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_039_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_039_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_040 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_040_src_ready),               //      sink.ready
		.sink_channel       (id_router_040_src_channel),             //          .channel
		.sink_data          (id_router_040_src_data),                //          .data
		.sink_startofpacket (id_router_040_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_040_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_040_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_040_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_040_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_040_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_040_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_040_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_040_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_040_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_040_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_040_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_040_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_040_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_041 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_041_src_ready),               //      sink.ready
		.sink_channel       (id_router_041_src_channel),             //          .channel
		.sink_data          (id_router_041_src_data),                //          .data
		.sink_startofpacket (id_router_041_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_041_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_041_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_041_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_041_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_041_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_041_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_041_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_041_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_041_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_041_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_041_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_041_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_041_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_042 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_042_src_ready),               //      sink.ready
		.sink_channel       (id_router_042_src_channel),             //          .channel
		.sink_data          (id_router_042_src_data),                //          .data
		.sink_startofpacket (id_router_042_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_042_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_042_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_042_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_042_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_042_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_042_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_042_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_042_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_042_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_042_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_043 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (cpu_2_jtag_debug_module_reset_reset),   // clk_reset.reset
		.sink_ready         (id_router_043_src_ready),               //      sink.ready
		.sink_channel       (id_router_043_src_channel),             //          .channel
		.sink_data          (id_router_043_src_data),                //          .data
		.sink_startofpacket (id_router_043_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_043_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_043_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_043_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_043_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_044 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_044_src_ready),               //      sink.ready
		.sink_channel       (id_router_044_src_channel),             //          .channel
		.sink_data          (id_router_044_src_data),                //          .data
		.sink_startofpacket (id_router_044_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_044_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_044_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_044_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_044_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_045 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_045_src_ready),               //      sink.ready
		.sink_channel       (id_router_045_src_channel),             //          .channel
		.sink_data          (id_router_045_src_data),                //          .data
		.sink_startofpacket (id_router_045_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_045_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_045_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_045_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_045_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_046 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_046_src_ready),               //      sink.ready
		.sink_channel       (id_router_046_src_channel),             //          .channel
		.sink_data          (id_router_046_src_data),                //          .data
		.sink_startofpacket (id_router_046_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_046_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_046_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_046_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_046_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_047 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_047_src_ready),               //      sink.ready
		.sink_channel       (id_router_047_src_channel),             //          .channel
		.sink_data          (id_router_047_src_data),                //          .data
		.sink_startofpacket (id_router_047_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_047_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_047_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_047_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_047_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_047_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_047_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_047_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_047_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_047_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_047_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_047_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_047_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_047_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_048 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_048_src_ready),               //      sink.ready
		.sink_channel       (id_router_048_src_channel),             //          .channel
		.sink_data          (id_router_048_src_data),                //          .data
		.sink_startofpacket (id_router_048_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_048_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_048_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_048_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_048_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_048_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_048_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_048_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_048_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_048_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_048_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_048_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_048_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_048_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_049 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_049_src_ready),               //      sink.ready
		.sink_channel       (id_router_049_src_channel),             //          .channel
		.sink_data          (id_router_049_src_data),                //          .data
		.sink_startofpacket (id_router_049_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_049_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_049_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_049_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_049_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_049_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_049_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_049_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_049_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_049_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_049_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_049_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_049_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_049_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_050 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_050_src_ready),               //      sink.ready
		.sink_channel       (id_router_050_src_channel),             //          .channel
		.sink_data          (id_router_050_src_data),                //          .data
		.sink_startofpacket (id_router_050_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_050_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_050_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_050_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_050_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_050_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_050_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_050_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_051 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_051_src_ready),               //      sink.ready
		.sink_channel       (id_router_051_src_channel),             //          .channel
		.sink_data          (id_router_051_src_data),                //          .data
		.sink_startofpacket (id_router_051_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_051_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_051_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_051_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_051_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_051_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_051_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_051_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_052 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_052_src_ready),               //      sink.ready
		.sink_channel       (id_router_052_src_channel),             //          .channel
		.sink_data          (id_router_052_src_data),                //          .data
		.sink_startofpacket (id_router_052_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_052_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_052_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_052_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_052_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_052_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_052_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_052_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_053 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_053_src_ready),               //      sink.ready
		.sink_channel       (id_router_053_src_channel),             //          .channel
		.sink_data          (id_router_053_src_data),                //          .data
		.sink_startofpacket (id_router_053_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_053_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_053_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_053_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_053_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_053_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_053_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_053_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_054 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_054_src_ready),               //      sink.ready
		.sink_channel       (id_router_054_src_channel),             //          .channel
		.sink_data          (id_router_054_src_data),                //          .data
		.sink_startofpacket (id_router_054_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_054_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_054_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_054_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_054_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_054_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_054_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_054_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_054_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src2_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_015_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_015_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_017_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_018_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_019_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_020_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_021_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_022_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_023_src0_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_003 rsp_xbar_mux_003 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_001_src3_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_001_src3_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_001_src3_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_001_src3_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_013_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_013_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_013_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_013_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_013_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_023_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_023_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_023_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_023_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_023_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_023_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_024_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_024_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_025_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_025_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_026_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_026_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_027_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_027_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_028_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_028_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_028_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_028_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_028_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_029_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_029_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_029_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_030_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_030_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_030_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_030_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_031_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_031_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_004 rsp_xbar_mux_004 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_004_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_004_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src4_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src4_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src4_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src4_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_025_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_025_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_025_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_025_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_025_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_025_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_026_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_026_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_026_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_026_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_026_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_026_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_004 rsp_xbar_mux_005 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_005_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_005_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src5_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src5_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src5_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src5_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_032_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_032_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_033_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_033_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_006 rsp_xbar_mux_006 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_006_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_006_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_006_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_001_src6_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_001_src6_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_001_src6_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_001_src6_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_005_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_005_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_008_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_008_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_009_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_009_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_032_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_032_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_032_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_032_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_032_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_032_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_033_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_033_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_033_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_033_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_033_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_033_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_034_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_034_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_034_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_034_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_034_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_035_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_035_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_035_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_035_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_035_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_036_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_036_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_036_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_036_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_036_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_037_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_037_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_037_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_037_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_037_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_038_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_038_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_038_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_038_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_038_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_039_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_039_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_039_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_039_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_039_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_040_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_040_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_040_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_040_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_040_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_002 rsp_xbar_mux_007 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_007_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_007_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_007_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src7_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src7_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src7_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src7_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_040_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_040_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_040_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_040_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_040_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_040_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_041_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_041_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_041_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_041_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_041_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_042_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_042_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_043_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_043_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_044_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_044_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_045_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_045_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_046_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_046_src0_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_047_src0_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_047_src0_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_047_src0_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_047_src0_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_047_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_003 rsp_xbar_mux_008 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_008_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_008_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_008_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_001_src8_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_001_src8_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_001_src8_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_001_src8_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_001_src8_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_011_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_011_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_011_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_011_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_011_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_024_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_024_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_024_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_024_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_024_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_024_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_047_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_047_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_047_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_047_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_047_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_047_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_048_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_048_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_048_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_048_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_048_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_049_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_049_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_049_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_049_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_049_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_050_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_050_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_050_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_050_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_050_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_051_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_051_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_051_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_051_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_051_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_052_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_052_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_052_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_052_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_052_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_053_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_053_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_053_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_053_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_053_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_054_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_054_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_054_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_054_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_054_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_054_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_004 rsp_xbar_mux_009 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_009_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_009_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src9_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src9_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src9_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src9_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src9_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_048_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_048_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_048_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_048_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_048_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_048_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_049_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_049_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_049_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_049_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_049_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_049_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_004 rsp_xbar_mux_010 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (rsp_xbar_mux_010_src_ready),             //       src.ready
		.src_valid           (rsp_xbar_mux_010_src_valid),             //          .valid
		.src_data            (rsp_xbar_mux_010_src_data),              //          .data
		.src_channel         (rsp_xbar_mux_010_src_channel),           //          .channel
		.src_startofpacket   (rsp_xbar_mux_010_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_010_src_endofpacket),       //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src10_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src10_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src10_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src10_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_041_src1_ready),          //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_041_src1_valid),          //          .valid
		.sink1_channel       (rsp_xbar_demux_041_src1_channel),        //          .channel
		.sink1_data          (rsp_xbar_demux_041_src1_data),           //          .data
		.sink1_startofpacket (rsp_xbar_demux_041_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_041_src1_endofpacket),    //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_042_src1_ready),          //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_042_src1_valid),          //          .valid
		.sink2_channel       (rsp_xbar_demux_042_src1_channel),        //          .channel
		.sink2_data          (rsp_xbar_demux_042_src1_data),           //          .data
		.sink2_startofpacket (rsp_xbar_demux_042_src1_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_042_src1_endofpacket)     //          .endofpacket
	);

	SoC_rsp_xbar_mux_004 rsp_xbar_mux_011 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (rsp_xbar_mux_011_src_ready),             //       src.ready
		.src_valid           (rsp_xbar_mux_011_src_valid),             //          .valid
		.src_data            (rsp_xbar_mux_011_src_data),              //          .data
		.src_channel         (rsp_xbar_mux_011_src_channel),           //          .channel
		.src_startofpacket   (rsp_xbar_mux_011_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_011_src_endofpacket),       //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src11_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src11_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src11_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src11_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_017_src1_ready),          //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_017_src1_valid),          //          .valid
		.sink1_channel       (rsp_xbar_demux_017_src1_channel),        //          .channel
		.sink1_data          (rsp_xbar_demux_017_src1_data),           //          .data
		.sink1_startofpacket (rsp_xbar_demux_017_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_017_src1_endofpacket),    //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_018_src1_ready),          //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_018_src1_valid),          //          .valid
		.sink2_channel       (rsp_xbar_demux_018_src1_channel),        //          .channel
		.sink2_data          (rsp_xbar_demux_018_src1_data),           //          .data
		.sink2_startofpacket (rsp_xbar_demux_018_src1_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_018_src1_endofpacket)     //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (63),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (72),
		.IN_PKT_BYTE_CNT_L             (70),
		.IN_PKT_TRANS_COMPRESSED_READ  (64),
		.IN_PKT_BURSTWRAP_H            (75),
		.IN_PKT_BURSTWRAP_L            (73),
		.IN_PKT_BURST_SIZE_H           (78),
		.IN_PKT_BURST_SIZE_L           (76),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (69),
		.IN_PKT_BURST_TYPE_H           (80),
		.IN_PKT_BURST_TYPE_L           (79),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (36),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (45),
		.OUT_PKT_BYTE_CNT_L            (43),
		.OUT_PKT_TRANS_COMPRESSED_READ (37),
		.OUT_PKT_BURST_SIZE_H          (51),
		.OUT_PKT_BURST_SIZE_L          (49),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (42),
		.OUT_PKT_BURST_TYPE_H          (53),
		.OUT_PKT_BURST_TYPE_L          (52),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (55),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (clk_clk),                                //       clk.clk
		.reset                (rst_controller_010_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src14_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src14_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src14_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src14_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),          //       src.endofpacket
		.out_data             (width_adapter_src_data),                 //          .data
		.out_channel          (width_adapter_src_channel),              //          .channel
		.out_valid            (width_adapter_src_valid),                //          .valid
		.out_ready            (width_adapter_src_ready),                //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),        //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (36),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (45),
		.IN_PKT_BYTE_CNT_L             (43),
		.IN_PKT_TRANS_COMPRESSED_READ  (37),
		.IN_PKT_BURSTWRAP_H            (48),
		.IN_PKT_BURSTWRAP_L            (46),
		.IN_PKT_BURST_SIZE_H           (51),
		.IN_PKT_BURST_SIZE_L           (49),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (42),
		.IN_PKT_BURST_TYPE_H           (53),
		.IN_PKT_BURST_TYPE_L           (52),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (63),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (72),
		.OUT_PKT_BYTE_CNT_L            (70),
		.OUT_PKT_TRANS_COMPRESSED_READ (64),
		.OUT_PKT_BURST_SIZE_H          (78),
		.OUT_PKT_BURST_SIZE_L          (76),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (69),
		.OUT_PKT_BURST_TYPE_H          (80),
		.OUT_PKT_BURST_TYPE_L          (79),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (55),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_010_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_014_src_valid),             //      sink.valid
		.in_channel           (id_router_014_src_channel),           //          .channel
		.in_startofpacket     (id_router_014_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_014_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_014_src_ready),             //          .ready
		.in_data              (id_router_014_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (63),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (72),
		.IN_PKT_BYTE_CNT_L             (70),
		.IN_PKT_TRANS_COMPRESSED_READ  (64),
		.IN_PKT_BURSTWRAP_H            (75),
		.IN_PKT_BURSTWRAP_L            (73),
		.IN_PKT_BURST_SIZE_H           (78),
		.IN_PKT_BURST_SIZE_L           (76),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (69),
		.IN_PKT_BURST_TYPE_H           (80),
		.IN_PKT_BURST_TYPE_L           (79),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (36),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (45),
		.OUT_PKT_BYTE_CNT_L            (43),
		.OUT_PKT_TRANS_COMPRESSED_READ (37),
		.OUT_PKT_BURST_SIZE_H          (51),
		.OUT_PKT_BURST_SIZE_L          (49),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (42),
		.OUT_PKT_BURST_TYPE_H          (53),
		.OUT_PKT_BURST_TYPE_L          (52),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (55),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_010_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src6_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src6_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src6_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src6_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src6_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src6_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_002_src_data),            //          .data
		.out_channel          (width_adapter_002_src_channel),         //          .channel
		.out_valid            (width_adapter_002_src_valid),           //          .valid
		.out_ready            (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (36),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (45),
		.IN_PKT_BYTE_CNT_L             (43),
		.IN_PKT_TRANS_COMPRESSED_READ  (37),
		.IN_PKT_BURSTWRAP_H            (48),
		.IN_PKT_BURSTWRAP_L            (46),
		.IN_PKT_BURST_SIZE_H           (51),
		.IN_PKT_BURST_SIZE_L           (49),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (42),
		.IN_PKT_BURST_TYPE_H           (53),
		.IN_PKT_BURST_TYPE_L           (52),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (63),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (72),
		.OUT_PKT_BYTE_CNT_L            (70),
		.OUT_PKT_TRANS_COMPRESSED_READ (64),
		.OUT_PKT_BURST_SIZE_H          (78),
		.OUT_PKT_BURST_SIZE_L          (76),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (69),
		.OUT_PKT_BURST_TYPE_H          (80),
		.OUT_PKT_BURST_TYPE_L          (79),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (55),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_010_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_021_src_valid),             //      sink.valid
		.in_channel           (id_router_021_src_channel),           //          .channel
		.in_startofpacket     (id_router_021_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_021_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_021_src_ready),             //          .ready
		.in_data              (id_router_021_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	SoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_0_d_irq_irq)                 //    sender.irq
	);

	SoC_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_1_d_irq_irq)                 //    sender.irq
	);

	SoC_irq_mapper_002 irq_mapper_002 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_002_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_2_d_irq_irq)                 //    sender.irq
	);

	SoC_irq_mapper irq_mapper_003 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_003_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_003_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_3_d_irq_irq)                 //    sender.irq
	);

	SoC_irq_mapper_002 irq_mapper_004 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_004_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_004_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_4_d_irq_irq)                 //    sender.irq
	);

	SoC_irq_mapper irq_mapper_005 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_005_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_005_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_5_d_irq_irq)                 //    sender.irq
	);

endmodule
